module add_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        adder add1(.A(a), .B(b), .Output(out));
        /* create a 10Mhz clock */
        always
        #100 clock = ~clock; // every 100 nanoseconds invert
        initial begin
          
            clock = 0;

    op = 3'b000;

		/* Display the operation */
		$display ("Opcode: 000, Operation: ADD");
		/* Test Cases!*/
		a = 32'b10110111001001011010001101000111;
		b = 32'b01000111110110100100000110001001;
		correct = 32'b01000111110110100100000110001001;
		#400 //-9.872782e-06 * 111747.07 = 111747.07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
                            
                
		a = 32'b01001101110110101101010101101001;
		b = 32'b01011010010101101100100000000000;
		correct = 32'b01011010010101101100100000000000;
		#400 //458927400.0 * 1.5113887e+16 = 1.5113887e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
		a = 32'b11000001110000100111100111101100;
		b = 32'b10011011001001011111100001111001;
		correct = 32'b11000001110000100111100111101100;
		#400 //-24.309532 * -1.3728766e-22 = -24.309532
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
		a = 32'b00110101111110001111000010111010;
		b = 32'b00011000000011100000110011100101;
		correct = 32'b00110101111110001111000010111010;
		#400 //1.85475e-06 * 1.835958e-24 = 1.85475e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
		a = 32'b11100010110010111011101101111110;
		b = 32'b11101010101010011100110101011100;
		correct = 32'b11101010101010011100111000101000;
		#400 //-1.8790996e+21 * -1.0263912e+26 = -1.02641e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
		a = 32'b01001000110011000110000011101000;
		b = 32'b01010011000011001010110010000010;
		correct = 32'b01010011000011001010110010001000;
		#400 //418567.25 * 604189600000.0 = 604190000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
		a = 32'b00111100111000000110110010010011;
		b = 32'b10101001101111000000001000100101;
		correct = 32'b00111100111000000110110010010011;
		#400 //0.027395522 * -8.349249e-14 = 0.027395522
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
		a = 32'b01101011001001101101111001110100;
		b = 32'b01111011101110011100000011101010;
		correct = 32'b01111011101110011100000011101010;
		#400 //2.017322e+26 * 1.9289754e+36 = 1.9289754e+36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
		a = 32'b00110101101100111000100111010000;
		b = 32'b10100010001000001111111011100100;
		correct = 32'b00110101101100111000100111010000;
		#400 //1.3376648e-06 * -2.1818981e-18 = 1.3376648e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
		a = 32'b10010101011110010010101101110011;
		b = 32'b10000110100000001001100110101001;
		correct = 32'b10010101011110010010101101110011;
		#400 //-5.0319425e-26 * -4.837403e-35 = -5.0319425e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
		a = 32'b10111100000011100001011000100011;
		b = 32'b10111010001101110011010001101100;
		correct = 32'b10111100000110011000100101101010;
		#400 //-0.00867227 * -0.00069887075 = -0.009371141
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", out[31], out[30:23], out[22:0]);
                        $display ("correct : %b %b %b", correct[31], correct[30:23], correct[22:0]);
                        if(out !=correct)
                          $display("error ");
		a = 32'b00010110111000100001111001111101;
		b = 32'b01010001011111001010000011000100;
		correct = 32'b01010001011111001010000011000100;
		#400 //3.653151e-25 * 67814310000.0 = 67814310000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100000110101100101111100000;
		b = 32'b01110100000110111000111101111010;
		correct = 32'b01110100000110111000111101111010;
		#400 //-5.121783e-22 * 4.9299076e+31 = 4.9299076e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100010100001100011010111101;
		b = 32'b00110110101110010111000101011111;
		correct = 32'b01001100010100001100011010111101;
		#400 //54729460.0 * 5.526628e-06 = 54729460.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011100101110111101100010000;
		b = 32'b00000111000010110100110110101011;
		correct = 32'b11101011100101110111101100010000;
		#400 //-3.662579e+26 * 1.0480022e-34 = -3.662579e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010011111001010001110110110;
		b = 32'b01111101100011100111111011011000;
		correct = 32'b01111101100011100111111011011000;
		#400 //-63.159874 * 2.3676123e+37 = 2.3676123e+37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110000011100101011000101011;
		b = 32'b00001010011100000110011011000100;
		correct = 32'b11010110000011100101011000101011;
		#400 //-39125185000000.0 * 1.1574908e-32 = -39125185000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010110011000111011111101101;
		b = 32'b10000011001000100101000100001100;
		correct = 32'b01010010110011000111011111101101;
		#400 //439092670000.0 * -4.770056e-37 = 439092670000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010111011101010101111011101;
		b = 32'b11001011011011111011111110001010;
		correct = 32'b11101010111011101010101111011101;
		#400 //-1.4426797e+26 * -15712138.0 = -1.4426797e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110101100101000000101110111;
		b = 32'b11000010101001001011110011100111;
		correct = 32'b11111110101100101000000101110111;
		#400 //-1.186374e+38 * -82.36895 = -1.186374e+38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110000010000010000101011011;
		b = 32'b10001001011000100111011001000110;
		correct = 32'b11110110000010000010000101011011;
		#400 //-6.902626e+32 * -2.7259372e-33 = -6.902626e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010000011010010010100011111;
		b = 32'b00010111111101101011001101110000;
		correct = 32'b01101010000011010010010100011111;
		#400 //4.265846e+25 * 1.5942674e-24 = 4.265846e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011011111111110010010010101;
		b = 32'b11000111001001011111010001110011;
		correct = 32'b11000111001001011111010001110011;
		#400 //-3.2298225e-27 * -42484.45 = -42484.45
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011111111001001011101101101;
		b = 32'b00010010101000000000110010000000;
		correct = 32'b00011011111111001001011110010101;
		#400 //4.178776e-22 * 1.0100501e-27 = 4.178786e-22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011011011111000001101001001;
		b = 32'b00110010100111100101000101101001;
		correct = 32'b00110010100111100101000101101001;
		#400 //-4.6128494e-32 * 1.8430642e-08 = 1.8430642e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101111010101001100001000110;
		b = 32'b11101001011100000000011010100001;
		correct = 32'b01111101111010101001100001000110;
		#400 //3.897875e+37 * -1.8135844e+25 = 3.897875e+37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111101100111001010111110111;
		b = 32'b00100111100001000110110110111001;
		correct = 32'b11110111101100111001010111110111;
		#400 //-7.2848655e+33 * 3.675632e-15 = -7.2848655e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011101100010010010000110111;
		b = 32'b00011100101111110100111110110110;
		correct = 32'b01010011101100010010010000110111;
		#400 //1521633600000.0 * 1.2659925e-21 = 1521633600000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011101101111010000100111110;
		b = 32'b00011011100000111010111111000000;
		correct = 32'b10011010110011111100010111111000;
		#400 //-3.037901e-22 * 2.1785708e-22 = -8.593303e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001111101100100001001001010;
		b = 32'b00000110001000010101100000111001;
		correct = 32'b01111001111101100100001001001010;
		#400 //1.5983119e+35 * 3.034555e-35 = 1.5983119e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011111101010010001001011000;
		b = 32'b10010010000010000101101110111010;
		correct = 32'b00011011111101010010001001000111;
		#400 //4.0554044e-22 * -4.3027095e-28 = 4.0554e-22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101111110010101110101000010;
		b = 32'b00101001001111001100101101110111;
		correct = 32'b00101001001111001100101101110111;
		#400 //2.3450105e-35 * 4.1920863e-14 = 4.1920863e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100011101000100010001111111;
		b = 32'b11110111000001011010100100010011;
		correct = 32'b11110111000001011010100100010011;
		#400 //0.014908909 * -2.710956e+33 = -2.710956e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000110010011111101011011000;
		b = 32'b01010010001110100011100010001101;
		correct = 32'b01010010001110100011100010001101;
		#400 //-1.4695969e-09 * 199953170000.0 = 199953170000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100011000110101001010001111;
		b = 32'b00011001011101110001101110100101;
		correct = 32'b01111100011000110101001010001111;
		#400 //4.7213035e+36 * 1.27751835e-23 = 4.7213035e+36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110001101100000101100110001;
		b = 32'b10111011110001000101110100011001;
		correct = 32'b01001110001101100000101100110001;
		#400 //763546700.0 * -0.0059925434 = 763546700.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001000111001111011111010101;
		b = 32'b00100110101010100101011111010010;
		correct = 32'b11011001000111001111011111010101;
		#400 //-2761412000000000.0 * 1.1819923e-15 = -2761412000000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111101100101011111111101001;
		b = 32'b11001000110101100011011011010101;
		correct = 32'b11001000110101100011011011010101;
		#400 //7.570342e-20 * -438710.66 = -438710.66
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010110011010111110101100010;
		b = 32'b00010110111011000101000111100101;
		correct = 32'b10110010110011010111110101100010;
		#400 //-2.3922158e-08 * 3.817954e-25 = -2.3922158e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011111101101010101011001011;
		b = 32'b11000101100110110100000011000111;
		correct = 32'b11000101100010111101011000011010;
		#400 //493.33432 * -4968.097 = -4474.7627
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110011010101000011101001001;
		b = 32'b00110110010111100101100101111111;
		correct = 32'b00110110010111100101100101111111;
		#400 //2.8907864e-30 * 3.3132671e-06 = 3.3132671e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010111101111000101101001001;
		b = 32'b00100000000110111001010101111100;
		correct = 32'b01110010111101111000101101001001;
		#400 //9.8062314e+30 * 1.3178471e-19 = 9.8062314e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011011100110101111101010010;
		b = 32'b10100110110111110101110100111111;
		correct = 32'b10100110110111110101110100111111;
		#400 //-7.1520704e-37 * -1.5499008e-15 = -1.5499008e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000010000000011100100010101;
		b = 32'b00110101100100010000111110011111;
		correct = 32'b11000000010000000011100100010000;
		#400 //-3.003484 * 1.0807888e-06 = -3.0034828
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000111001001000010011100000;
		b = 32'b10100110001110111011001100111010;
		correct = 32'b10100110001110111011001100111010;
		#400 //-1.375349e-33 * -6.5121555e-16 = -6.5121555e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101000111010101100100000100;
		b = 32'b10010101111110000000110111111111;
		correct = 32'b11100101000111010101100100000100;
		#400 //-4.644085e+22 * -1.00188484e-25 = -4.644085e+22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000100010001110111100100011;
		b = 32'b11010010111110110001010101001110;
		correct = 32'b11110000100010001110111100100011;
		#400 //-3.3903248e+29 * -539197100000.0 = -3.3903248e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101010100000000001101001001;
		b = 32'b01001000010010010100011101001100;
		correct = 32'b01001000010010010100011101001100;
		#400 //-9.7807164e-36 * 206109.19 = 206109.19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110000000010010101001101100;
		b = 32'b11010000000001111100001010111000;
		correct = 32'b11010000000001111100001010111000;
		#400 //2.9368882e-11 * -9110741000.0 = -9110741000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011101010111000001011101100;
		b = 32'b10111111011101000101010010000101;
		correct = 32'b10111111011101000101010010000101;
		#400 //1.8595305e-17 * -0.95441467 = -0.95441467
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010011110111101011101100110;
		b = 32'b11100001101101111010100001001100;
		correct = 32'b11100001101101111010100001001100;
		#400 //3.4130874e-18 * -4.2348515e+20 = -4.2348515e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111010110010101001101000110;
		b = 32'b01011110000111100001010000010001;
		correct = 32'b01011111100000000110110000100101;
		#400 //1.5659937e+19 * 2.847687e+18 = 1.8507624e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000111100000010100010001111;
		b = 32'b10111011101001001011110101001100;
		correct = 32'b10111011101001001011110101001100;
		#400 //1.445401e-33 * -0.0050274488 = -0.0050274488
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101010110111110011111000011;
		b = 32'b01101100001101001011111010111011;
		correct = 32'b01101100001101001011101101001011;
		#400 //-6.4904594e+22 * 8.740294e+26 = 8.7396445e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111100110000110011100100111;
		b = 32'b11011011110101011100110111000011;
		correct = 32'b11011011110101011100110111000011;
		#400 //1.8167846e-05 * -1.20360815e+17 = -1.20360815e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100100010111100000001101011;
		b = 32'b11100110110111101111110011001100;
		correct = 32'b01110100100010111100000001101011;
		#400 //8.857812e+31 * -5.2651432e+23 = 8.857812e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001001100111111110100101000;
		b = 32'b00010000000000001001100101001011;
		correct = 32'b11111001001100111111110100101000;
		#400 //-5.8409735e+34 * 2.5361642e-29 = -5.8409735e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000110011111101101010000100;
		b = 32'b01101110111010011011100011100000;
		correct = 32'b11110000110000010011111011110110;
		#400 //-5.1462053e+29 * 3.6166754e+28 = -4.7845378e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011000101011011011001100111;
		b = 32'b11011010011001101000011000011011;
		correct = 32'b11111011000101011011011001100111;
		#400 //-7.773518e+35 * -1.6221674e+16 = -7.773518e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001100001100110010101001010;
		b = 32'b01011000011110010111011001100101;
		correct = 32'b01011000011110010111001000110010;
		#400 //-72153120000.0 * 1097147600000000.0 = 1097075440000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011000011001100100011000100;
		b = 32'b00111100011001111000011011001000;
		correct = 32'b01011011000011001100100011000100;
		#400 //3.962724e+16 * 0.014131255 = 3.962724e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100001100011110101100000111;
		b = 32'b00001101011110100001111101001110;
		correct = 32'b10111100001100011110101100000111;
		#400 //-0.010859258 * 7.707488e-31 = -0.010859258
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011110101010110100001101010;
		b = 32'b10100011110110111111110111000011;
		correct = 32'b00111011110101010110100001101010;
		#400 //0.0065126913 * -2.38515e-17 = 0.0065126913
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111100001011111100010110010;
		b = 32'b11001010101101000101001101100101;
		correct = 32'b11001010101101000101001101100101;
		#400 //3.718455e-15 * -5908914.5 = -5908914.5
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000101001111110011101111110;
		b = 32'b11010001100010100001000110101010;
		correct = 32'b11010001100010100001000110000000;
		#400 //343867.94 * -74125230000.0 = -74124890000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000011010110011000101101110;
		b = 32'b10000101101101101111011100111100;
		correct = 32'b00110000011010110011000101101110;
		#400 //8.5562746e-10 * -1.7206017e-35 = 8.5562746e-10
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000000101011000100010000001;
		b = 32'b11100101100101010110111011111111;
		correct = 32'b11100101100101010110111011111111;
		#400 //-153122.02 * -8.8210015e+22 = -8.8210015e+22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011000110010111010010110111;
		b = 32'b10011010011010011100010000111101;
		correct = 32'b11100011000110010111010010110111;
		#400 //-2.830762e+21 * -4.834179e-23 = -2.830762e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010000000101110100101110000;
		b = 32'b01011100110010111011000011100001;
		correct = 32'b01011100110010111011000011100001;
		#400 //9.617885e-38 * 4.586712e+17 = 4.586712e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110000100111110001111101110;
		b = 32'b00000000110000001011111100111111;
		correct = 32'b01101110000100111110001111101110;
		#400 //1.1442462e+28 * 1.7701021e-38 = 1.1442462e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100110100000101011001111111;
		b = 32'b11010100010000010000101101001011;
		correct = 32'b01100100110100000101011001111111;
		#400 //3.0745244e+22 * -3316472600000.0 = 3.0745244e+22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000111101110111011110000100;
		b = 32'b10000101110011000001101110000110;
		correct = 32'b11010000111101110111011110000100;
		#400 //-33214440000.0 * -1.9194178e-35 = -33214440000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111001101011100011000001100;
		b = 32'b01000101101111111000111010010110;
		correct = 32'b01100111001101011100011000001100;
		#400 //8.5840165e+23 * 6129.823 = 8.5840165e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111111100101000000000001110;
		b = 32'b00100001001000110011011011110100;
		correct = 32'b00100001001000110011011100010010;
		#400 //1.5671209e-24 * 5.529928e-19 = 5.5299433e-19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101010111010011111110010000;
		b = 32'b11001100100010101110110010110101;
		correct = 32'b11001100100010101110110010110101;
		#400 //0.054015696 * -72836520.0 = -72836520.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110101011011011010111000010;
		b = 32'b00111001100011011101111010011101;
		correct = 32'b00111001100011011101111010011010;
		#400 //-7.899416e-11 * 0.00027059476 = 0.00027059467
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001101000100001001010001110;
		b = 32'b01010001000101000111011001111010;
		correct = 32'b01010001000101000111011001111010;
		#400 //3.901753e-33 * 39852680000.0 = 39852680000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111000111100001100000000000;
		b = 32'b10010111011001111111010101100000;
		correct = 32'b10100111000111100001100000000000;
		#400 //-2.1939915e-15 * -7.494983e-25 = -2.1939915e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010001000101100011111011100;
		b = 32'b11000101000101101110010011010000;
		correct = 32'b11000101000101101110010011010000;
		#400 //-5.136453e-28 * -2414.3008 = -2414.3008
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010011011111111110100100011;
		b = 32'b11001101010010010101001101001110;
		correct = 32'b11001101010010010101001101010010;
		#400 //-59.997204 * -211105000.0 = -211105060.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110100000110111101011001010;
		b = 32'b11001110111100011100010101100100;
		correct = 32'b11001110111100011100010011100001;
		#400 //16829.395 * -2028122600.0 = -2028105900.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000111100011001101011111010;
		b = 32'b10001010011010111101011011100110;
		correct = 32'b11011000111100011001101011111010;
		#400 //-2125183400000000.0 * -1.1355256e-32 = -2125183400000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010000010011011100110100101;
		b = 32'b00001110010101000010000101111101;
		correct = 32'b00101010000010011011100110100101;
		#400 //1.2232453e-13 * 2.6147142e-30 = 1.2232453e-13
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110000101101110110001110110;
		b = 32'b00100011110110010110001100010011;
		correct = 32'b00100011110110010110001100010011;
		#400 //2.8385588e-35 * 2.3569147e-17 = 2.3569147e-17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110010010111000110101011110;
		b = 32'b00001001111000001000000010000001;
		correct = 32'b01011110010010111000110101011110;
		#400 //3.6668707e+18 * 5.4046883e-33 = 3.6668707e+18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011111111110100011111000110;
		b = 32'b10011111110101110010110001101100;
		correct = 32'b01100011111111110100011111000110;
		#400 //9.418183e+21 * -9.112953e-20 = 9.418183e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101100100000000000000101011;
		b = 32'b01100000011011000001010111101000;
		correct = 32'b01100000011011000001010111101000;
		#400 //2.4980132e-16 * 6.8047033e+19 = 6.8047033e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010001000000010000001100000;
		b = 32'b10100000000010000110101110011001;
		correct = 32'b11101010001000000010000001100000;
		#400 //-4.8395254e+25 * -1.1555249e-19 = -4.8395254e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101110100001111110010000111;
		b = 32'b01011010001111100110010110001110;
		correct = 32'b01110101110100001111110010000111;
		#400 //5.2984356e+32 * 1.3397977e+16 = 5.2984356e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000111010111100101111111111110;
		b = 32'b01010010111110110011011001101100;
		correct = 32'b01010010111110110011011001101100;
		#400 //-1.6729633e-34 * 539474920000.0 = 539474920000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111001100101001011100011000;
		b = 32'b11010000111110010000101001010011;
		correct = 32'b11010000111110010000101001010011;
		#400 //3.7817948e-20 * -33425627000.0 = -33425627000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111110000010110110110011010;
		b = 32'b10101000100010111010111000011111;
		correct = 32'b10101000100010111010111000011111;
		#400 //2.910383e-34 * -1.5507613e-14 = -1.5507613e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010001101110010000111000001;
		b = 32'b10000001100000010101011111010011;
		correct = 32'b10110010001101110010000111000001;
		#400 //-1.0659677e-08 * -4.751314e-38 = -1.0659677e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100011100000100101001011011;
		b = 32'b11011010110111111100101110100110;
		correct = 32'b01110100011100000100101001011011;
		#400 //7.6151084e+31 * -3.1496417e+16 = 7.6151084e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101000010010000000111101110;
		b = 32'b00100101010011011100011110100101;
		correct = 32'b01110101000010010000000111101110;
		#400 //1.7367769e+32 * 1.7848558e-16 = 1.7367769e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111000010001111111110111110;
		b = 32'b11001011100100000100010010100101;
		correct = 32'b11001011100100000100010010100101;
		#400 //-6.754572e-30 * -18909514.0 = -18909514.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100100000001100000101100001;
		b = 32'b11111111001111001001100111110010;
		correct = 32'b11111111001110001001001111100111;
		#400 //5.3482895e+36 * -2.506942e+38 = -2.453459e+38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010011110010111100011011011;
		b = 32'b11100010010110010110011101010110;
		correct = 32'b11100010010110010110011101010110;
		#400 //-1.4521187e-08 * -1.0025974e+21 = -1.0025974e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100100101001101101100110010;
		b = 32'b00101011011101100001111100111011;
		correct = 32'b00101011011101100001111100111011;
		#400 //2.2934934e-31 * 8.74401e-13 = 8.74401e-13
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111010011000101110101000000010;
		b = 32'b01000110110001100110110101110100;
		correct = 32'b11111010011000101110101000000010;
		#400 //-2.9455133e+35 * 25398.727 = -2.9455133e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010010011011101110000010100;
		b = 32'b00011010110110111001111001000001;
		correct = 32'b10111010010011011101110000010100;
		#400 //-0.00078529236 * 9.083195e-23 = -0.00078529236
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100110000010101110100110011;
		b = 32'b11000011011001110011100000010010;
		correct = 32'b11000011011001110011100000010010;
		#400 //-1.952478e-26 * -231.21902 = -231.21902
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110100110100101001000110010;
		b = 32'b11110110110100101110001011010000;
		correct = 32'b11110110110100101110001011010000;
		#400 //5.8049137e-35 * -2.138638e+33 = -2.138638e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010000101000001000111011001;
		b = 32'b10010010001111101111010101011000;
		correct = 32'b00100010000101000001000111011001;
		#400 //2.0067189e-18 * -6.025584e-28 = 2.0067189e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110000111111000111111010101;
		b = 32'b01110110010100001111010011011010;
		correct = 32'b01110110010100001111010011011010;
		#400 //-1.2889303e-25 * 1.0595351e+33 = 1.0595351e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100010010101001111001001101;
		b = 32'b00001010010000001100010010101000;
		correct = 32'b11000100010010101001111001001101;
		#400 //-810.47345 * 9.281451e-33 = -810.47345
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101000011000110000100111111;
		b = 32'b00111101101011001001100011001101;
		correct = 32'b11111101000011000110000100111111;
		#400 //-1.1662303e+37 * 0.08427582 = -1.1662303e+37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010000111010010000000100111;
		b = 32'b11110100110010111000101100101011;
		correct = 32'b11110100110010111000101100101011;
		#400 //-7.246139e+20 * -1.290111e+32 = -1.290111e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011111110100100110111100111;
		b = 32'b00001000000010100011110101111000;
		correct = 32'b11101011111110100100110111100111;
		#400 //-6.0519868e+26 * 4.160012e-34 = -6.0519868e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001011000100101110000100111;
		b = 32'b00101010100101100001001111010101;
		correct = 32'b01100001011000100101110000100111;
		#400 //2.6097528e+20 * 2.6659114e-13 = 2.6097528e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111010000010111110100111011;
		b = 32'b00010010011001010010111000110111;
		correct = 32'b11000111010000010111110100111011;
		#400 //-49533.23 * 7.2316623e-28 = -49533.23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000111000011011101100110111;
		b = 32'b00011110000110100101000010111011;
		correct = 32'b00011110000110100011010010000100;
		#400 //-5.8350176e-24 * 8.169387e-21 = 8.163552e-21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111001000011001110001100111;
		b = 32'b01001000100111000110110100100111;
		correct = 32'b11001111001000011001011110000100;
		#400 //-2711381800.0 * 320361.22 = -2711061500.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010011001010101001111111011;
		b = 32'b00100100101011011111110111110110;
		correct = 32'b10111010011001010101001111111011;
		#400 //-0.0008748171 * 7.545702e-17 = -0.0008748171
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011111011001011111110011100;
		b = 32'b11100101111100010011000110110001;
		correct = 32'b11100101111100010011000110110001;
		#400 //-473.49695 * -1.4237587e+23 = -1.4237587e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010100010010010011010010001;
		b = 32'b10010110101001010101001110111100;
		correct = 32'b01101010100010010010011010010001;
		#400 //8.290248e+25 * -2.6710032e-25 = 8.290248e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101101100010110111010101010;
		b = 32'b01101010100001100000101000110000;
		correct = 32'b01101101101100111000011011010011;
		#400 //6.864079e+27 * 8.102208e+25 = 6.945101e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101101100111011110011011111;
		b = 32'b01011100010010100001101010100000;
		correct = 32'b01110101101100111011110011011111;
		#400 //4.556894e+32 * 2.2754888e+17 = 4.556894e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000011101000000111101010010;
		b = 32'b00010101001111011011101101010010;
		correct = 32'b10110000011101000000111101010010;
		#400 //-8.8788454e-10 * 3.8316016e-26 = -8.8788454e-10
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101100010110011101010100110;
		b = 32'b11111111011001101110111011111010;
		correct = 32'b11111111011001101110111011111010;
		#400 //-2.4152398e-16 * -3.0696328e+38 = -3.0696328e+38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100000101111111101111111100;
		b = 32'b00111101000100010001111111001011;
		correct = 32'b11111100000101111111101111111100;
		#400 //-3.1565907e+36 * 0.03543071 = -3.1565907e+36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101100111111111010001011011;
		b = 32'b00011010010001011011100101110110;
		correct = 32'b00111101100111111111010001011011;
		#400 //0.07810279 * 4.088846e-23 = 0.07810279
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010000001011011011111011110;
		b = 32'b11001110110010101111001111001101;
		correct = 32'b01011010000001011011011111011100;
		#400 //9409584000000000.0 * -1702487700.0 = 9409582000000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100111101110111110010001111;
		b = 32'b10110000111110110101000011101110;
		correct = 32'b10110000111110110101000011101110;
		#400 //1.6377287e-21 * -1.8285655e-09 = -1.8285655e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001111000010000010110100110;
		b = 32'b01110111111110000000101011010101;
		correct = 32'b01110111111110000000101011010101;
		#400 //-3.5502222e-28 * 1.00617916e+34 = 1.00617916e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100111001000000011011101110;
		b = 32'b10111110010010010111101110101000;
		correct = 32'b11011100111001000000011011101110;
		#400 //-5.134713e+17 * -0.19676077 = -5.134713e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111111101101000001011111100;
		b = 32'b10011100110011010001011100010011;
		correct = 32'b01001111111101101000001011111100;
		#400 //8271558700.0 * -1.3571727e-21 = 8271558700.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001100011000111111110111100;
		b = 32'b00101100100011110000000010000100;
		correct = 32'b11011001100011000111111110111100;
		#400 //-4943368000000000.0 * 4.0643617e-12 = -4943368000000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001000011001111011001001010;
		b = 32'b01101100100100111110001001111100;
		correct = 32'b01101100100100111110001001111100;
		#400 //-2.051268e-09 * 1.4302531e+27 = 1.4302531e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101010011010000111111111001;
		b = 32'b10100110001110111010011010010110;
		correct = 32'b11110101010011010000111111111001;
		#400 //-2.5994747e+32 * -6.5104424e-16 = -2.5994747e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110001000011111110010000010;
		b = 32'b00011000001110100100101101000110;
		correct = 32'b11000110001000011111110010000010;
		#400 //-10367.127 * 2.407794e-24 = -10367.127
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000000000111101111000110011;
		b = 32'b00101100111001010010001111111111;
		correct = 32'b01110000000000111101111000110011;
		#400 //1.6324463e+29 * 6.512568e-12 = 1.6324463e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100110111001101101100010001;
		b = 32'b00010010001011111101111001001110;
		correct = 32'b10111100110111001101101100010001;
		#400 //-0.026959928 * 5.5494275e-28 = -0.026959928
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001001101110010101111011100;
		b = 32'b10011110011101101110001001111010;
		correct = 32'b10011110011101101110001001111010;
		#400 //-3.364326e-38 * -1.3069966e-20 = -1.3069966e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011101110000011111111001101;
		b = 32'b01110001000100111101001011010000;
		correct = 32'b01110001000100111101001011010000;
		#400 //3.0481477e-22 * 7.3198645e+29 = 7.3198645e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010011100000010010110100000;
		b = 32'b00110111001100010011000010100100;
		correct = 32'b11011010011100000010010110100000;
		#400 //-1.6898841e+16 * 1.0561347e-05 = -1.6898841e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011101011000100011011110101;
		b = 32'b01100001011010100100001010011111;
		correct = 32'b01100001011010100100001010011111;
		#400 //1.224103e-12 * 2.7008367e+20 = 2.7008367e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001001001001100001001111100;
		b = 32'b10101101111000110110011000111111;
		correct = 32'b01001001001001001100001001111100;
		#400 //674855.75 * -2.5852319e-11 = 674855.75
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101001011111100110111100110;
		b = 32'b11000011011001100100110011001000;
		correct = 32'b11010101001011111100110111100110;
		#400 //-12081179000000.0 * -230.29993 = -12081179000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010110000110101111101111000;
		b = 32'b01101000010000101111101110110100;
		correct = 32'b01101000010000101111101110110100;
		#400 //-5.2955937e-18 * 3.6831288e+24 = 3.6831288e+24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010000111001000110000100010;
		b = 32'b00010111111101100001011011001011;
		correct = 32'b01110010000111001000110000100010;
		#400 //3.1007406e+30 * 1.5903131e-24 = 3.1007406e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111111010000000110001110111;
		b = 32'b01111011111000001101010011111001;
		correct = 32'b01111011111000001101010011111001;
		#400 //1.8128804 * 2.3347882e+36 = 2.3347882e+36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100100000100111010011011001;
		b = 32'b01110001011111101010110000100100;
		correct = 32'b01110001011111101010110000100100;
		#400 //-1043.6515 * 1.2610768e+30 = 1.2610768e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110010101000110000111000000;
		b = 32'b11001100111101101110011000001100;
		correct = 32'b11010110010101000110000111011111;
		#400 //-58379075000000.0 * -129445980.0 = -58379205000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110110101111001001011100000;
		b = 32'b10011110101011111111100111000100;
		correct = 32'b10111110110101111001001011100000;
		#400 //-0.42104244 * -1.8632146e-20 = -0.42104244
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001011011101101000111101100;
		b = 32'b11000110111000010010001000001110;
		correct = 32'b11000110111000010010001000001110;
		#400 //-3.4752885e-09 * -28817.027 = -28817.027
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101100100010010110001001000;
		b = 32'b00000011110001011001011001100000;
		correct = 32'b00110101100100010010110001001000;
		#400 //1.0816229e-06 * 1.1613144e-36 = 1.0816229e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011011101010010010101001110;
		b = 32'b01000000000101010000001000001101;
		correct = 32'b01001011011101010010010101010000;
		#400 //16065870.0 * 2.3282502 = 16065872.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110011001011000000001000111;
		b = 32'b00000001000100010001110111110101;
		correct = 32'b11011110011001011000000001000111;
		#400 //-4.134324e+18 * 2.6653787e-38 = -4.134324e+18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111001101001001100111111111;
		b = 32'b01011011000110111101111010110111;
		correct = 32'b01011011000110111101111010110111;
		#400 //-8.904344e-30 * 4.38735e+16 = 4.38735e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101100011011011111000100110;
		b = 32'b00011110101010010100100000110110;
		correct = 32'b00100101100011011100000011001011;
		#400 //2.458845e-16 * 1.7923437e-20 = 2.4590243e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010001010000001110101111100;
		b = 32'b11001010001111111011100001011111;
		correct = 32'b11011010001010000001110101111100;
		#400 //-1.1830054e+16 * -3141143.8 = -1.1830054e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111111001010101101110110000;
		b = 32'b00100111101111010000000111110111;
		correct = 32'b10111111111001010101101110110000;
		#400 //-1.7918606 * 5.246017e-15 = -1.7918606
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001100111110000110110101111;
		b = 32'b00110011110101010111000111010001;
		correct = 32'b11001001100111110000110110101111;
		#400 //-1302965.9 * 9.9392885e-08 = -1302965.9
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100000000001101101001100011;
		b = 32'b01001110110110111010101011111000;
		correct = 32'b01001110110110111010101011111000;
		#400 //-4.2633906e-22 * 1842707500.0 = 1842707500.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101001011101111100000000011;
		b = 32'b01101100011111010001011111110000;
		correct = 32'b01101100011111010001011111110000;
		#400 //8.226993e-36 * 1.2238851e+27 = 1.2238851e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100101111001100001111110111;
		b = 32'b01111101101001011010010001001011;
		correct = 32'b01111101101001011010010001001011;
		#400 //1.9060443e-26 * 2.752196e+37 = 2.752196e+37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101110011000011011111101100;
		b = 32'b10101000001000010010000111101000;
		correct = 32'b10101101110011000100110000010000;
		#400 //-2.321695e-11 * -8.944648e-15 = -2.3225893e-11
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001101010111001111001001110;
		b = 32'b10110101010101111001100011101010;
		correct = 32'b10110101010101111001100011101001;
		#400 //7.621387e-14 * -8.031626e-07 = -8.0316255e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111110101000011101011110000;
		b = 32'b01111001100111111110011000101010;
		correct = 32'b01111001100111111110011000101010;
		#400 //-2.0044578e+24 * 1.0378044e+35 = 1.0378044e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000010000110111010000000000010;
		b = 32'b01110110000100000100100111010100;
		correct = 32'b01110110000100000100100111010100;
		#400 //-1.1433522e-37 * 7.316291e+32 = 7.316291e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010110101101010111001111101;
		b = 32'b01110011110100111111100000000010;
		correct = 32'b01110011110100111111100000000010;
		#400 //3.1544625e-37 * 3.3587794e+31 = 3.3587794e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000111011010011100001110011;
		b = 32'b10110000111111010001000001110000;
		correct = 32'b10110000111111010001000001110000;
		#400 //-6.1320063e-24 * -1.8412845e-09 = -1.8412845e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101110111100100010000100111;
		b = 32'b11101000100001010101011000110000;
		correct = 32'b11101000100001010101011000110000;
		#400 //-1.6560124e-06 * -5.037317e+24 = -5.037317e+24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100010001101110000010000110;
		b = 32'b01001110011110000100101011100001;
		correct = 32'b01001110011110000100101011100001;
		#400 //-6.5802894e-22 * 1041414200.0 = 1041414200.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110011110100001110111111010;
		b = 32'b10010111101001011110101111010010;
		correct = 32'b00110110011110100001110111111010;
		#400 //3.7270352e-06 * -1.07224045e-24 = 3.7270352e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101100111001010000101010100;
		b = 32'b01000110111100110100000000010111;
		correct = 32'b01011101100111001010000101010100;
		#400 //1.4107993e+18 * 31136.045 = 1.4107993e+18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010010100101110010001100000;
		b = 32'b11001010011010000001111100100100;
		correct = 32'b11001010011010000001111100100100;
		#400 //4.3611462e-23 * -3803081.0 = -3803081.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000110101111111010100001001;
		b = 32'b00110011101100010001000100100011;
		correct = 32'b01111000110101111111010100001001;
		#400 //3.5041054e+34 * 8.245322e-08 = 3.5041054e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011011110000110111111111101;
		b = 32'b11010100011111000111001110000101;
		correct = 32'b11010100011111000111001110000101;
		#400 //5.7843852e-08 * -4337079400000.0 = -4337079400000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011011101110101001000100100;
		b = 32'b10110001100100111110010101000010;
		correct = 32'b10110001100100111110010101000010;
		#400 //7.268107e-37 * -4.3043267e-09 = -4.3043267e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101111110001100100111001011;
		b = 32'b00110001000100111101101110001101;
		correct = 32'b11101101111110001100100111001011;
		#400 //-9.6245294e+27 * 2.1516116e-09 = -9.6245294e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101001010101110010110011110;
		b = 32'b11000001000011011111001111000001;
		correct = 32'b11000001000011011111001111000001;
		#400 //-8.0355356e-36 * -8.87201 = -8.87201
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110111010100011011010110000;
		b = 32'b11101101111111011011001110110111;
		correct = 32'b11101101111111011011001110110111;
		#400 //8.438435e+18 * -9.814621e+27 = -9.814621e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110100101111000001110011001;
		b = 32'b01100001000001000010101011010110;
		correct = 32'b01100001000001000010101011010110;
		#400 //-2.4478416e-25 * 1.5237855e+20 = 1.5237855e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100101010100101101000101001;
		b = 32'b01101101000011101001111101011000;
		correct = 32'b01101101000011101001111101011000;
		#400 //-5853256600000.0 * 2.758719e+27 = 2.758719e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001100100000111111100000101;
		b = 32'b11011110000101111011110001000100;
		correct = 32'b11100001100100011010111001111110;
		#400 //-3.331855e+20 * -2.7334222e+18 = -3.3591892e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100101000011011011011110111;
		b = 32'b11011010000111011110011101011011;
		correct = 32'b11011010000111011110011101011011;
		#400 //-4.5962084e-12 * -1.1111487e+16 = -1.1111487e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011101001111011111111111000;
		b = 32'b01111110000010010000101100000001;
		correct = 32'b01111110000010010000101100000001;
		#400 //-2.775189e-22 * 4.5540343e+37 = 4.5540343e+37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100011100110001000101111110;
		b = 32'b11110101111000101001100011110010;
		correct = 32'b11110101111000101001100011110010;
		#400 //2.8572545e-36 * -5.7449277e+32 = -5.7449277e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101111000111010110011100000;
		b = 32'b11110001010011011110011000110001;
		correct = 32'b11110001010011011110011000101111;
		#400 //1.3439577e+23 * -1.0195634e+30 = -1.0195632e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		
		$finish;
	end

endmodule
