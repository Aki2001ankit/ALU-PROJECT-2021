`include "alu.v"


    module and_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .A(a),
                .B(b),
                .OpCode(op),
                .O(out)
            );
        /* create a 10Mhz clock */
        always
        #100 clock = ~clock; // every 100 nanoseconds invert
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, a, b, op, out);
            clock = 0;

    op = 3'b100;

		/* Display the operation */
		$display ("Opcode: 100, Operation: AND");
		/* Test Cases!*/
		a = 32'b01110010110010001000000001010001;
		b = 32'b01001110001010001000000100001000;
		correct = 32'b01000010000010001000000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110010111001001110000101000;
		b = 32'b00100011001111101110111011010000;
		correct = 32'b00100010000111001000110000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101010101000110111010000000;
		b = 32'b11101101100001010101110100010000;
		correct = 32'b11100101000001000100110000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010010001100001000011000000;
		b = 32'b10011101001110011011000001000100;
		correct = 32'b10001000000000000001000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100010101100100011110111101;
		b = 32'b00111001110100001010100100101101;
		correct = 32'b00010000010100000000000100101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000001100011101110000111001;
		b = 32'b10100001010100010110011010011101;
		correct = 32'b00000000000100010100010000011001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010101000111100100100000011;
		b = 32'b01111111110000110010111100011111;
		correct = 32'b01100010100000110000100100000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001101101011111000010001010;
		b = 32'b00111011110101001011110000100111;
		correct = 32'b00001001100101001011000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110110110110111011100101100;
		b = 32'b10111010101001111001010011010000;
		correct = 32'b00011010100000110001010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100000110010011100011100100;
		b = 32'b10110111010111011100100011101001;
		correct = 32'b10010100000110010000100011100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101001000110011001010011111;
		b = 32'b11100000011101001101101000010111;
		correct = 32'b01100000001000000001001000010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110011110011000001100100000;
		b = 32'b11000110010011010010011101100101;
		correct = 32'b00000110010010010000001100100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100001001001011000110101111;
		b = 32'b10111011001100111010000000100011;
		correct = 32'b10010000001000001010000000100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111001001101101100000000111;
		b = 32'b10001010101010001011100101111001;
		correct = 32'b10001010001000001001100000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110010100000100001101101101;
		b = 32'b01000010110110010010100011011101;
		correct = 32'b01000010010100000000000001001101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101110100011111100011101101;
		b = 32'b01011110101111010011001000100011;
		correct = 32'b01011100100100010011000000100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011110110111000110110001100;
		b = 32'b01011011101100111011101010110101;
		correct = 32'b00000011100100111000100010000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101000001101010001011010101;
		b = 32'b10111110101100110010010011010101;
		correct = 32'b00111100000000100010000011010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111010110110000111001000100;
		b = 32'b01100100100011100011011110100110;
		correct = 32'b01100100000010100000011000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111100010000110000110101001;
		b = 32'b11010010100101000001101001001011;
		correct = 32'b01000010100000000000000000001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110001000101110100010000000;
		b = 32'b00101010010101000000111101111101;
		correct = 32'b00101010000000000000100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110101111100000100110001101;
		b = 32'b11001100010110101000010000011101;
		correct = 32'b00000100000110100000000000001101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011100001001111010110100111;
		b = 32'b00010010110100111000110110111111;
		correct = 32'b00010010100000001000010110100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001101101110110110101001011001;
		b = 32'b11010110111111110101111111001101;
		correct = 32'b00000100101110110100101001001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011000000100001011100111001;
		b = 32'b11011101011110110010111100101001;
		correct = 32'b10001001000000100000011100101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101010100111011101011101110;
		b = 32'b01011100101101001011100101111001;
		correct = 32'b01001100000100001011100001101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100010110011000011101000000;
		b = 32'b00100010011001010001100110111100;
		correct = 32'b00100000010000010000000100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100101111100000110110000010;
		b = 32'b11000111110101000110100011101011;
		correct = 32'b11000100100101000000100010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000000100111000111000111010;
		b = 32'b11100101101100011100110000100010;
		correct = 32'b11100000000100011000110000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001011100011010110000010110;
		b = 32'b10100000011001110111011011100010;
		correct = 32'b10100000011000010010010000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110011100000111000010001110;
		b = 32'b01100101001100001110000111111101;
		correct = 32'b00100100001100000110000010001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111000110101010011101010100;
		b = 32'b10011011011101111010000001110100;
		correct = 32'b00000011000100101010000001010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010000001100010000110111111;
		b = 32'b00010111111001011110101110011011;
		correct = 32'b00010010000001000010000110011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111100110011000001101011101;
		b = 32'b01001000011101011011100001001010;
		correct = 32'b00001000000100011000000001001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001100010110100101000000001;
		b = 32'b01010010000100000011001000110100;
		correct = 32'b01010000000000000000001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101101101001001111101100010;
		b = 32'b00110010000000001000110110110110;
		correct = 32'b00110000000000001000110100100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011101011011100001010101010;
		b = 32'b00100000010000101001101101100101;
		correct = 32'b00100000000000001000001000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011101001000010011100000010;
		b = 32'b11000100010011000001101101110001;
		correct = 32'b11000000000001000000001100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010111001110101001001010011;
		b = 32'b00000101101000011010111011010100;
		correct = 32'b00000000101000010000001001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011001000111101111110011110;
		b = 32'b01100111011100000111111111110000;
		correct = 32'b01100011001000000101111110010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100111011111010111000001111;
		b = 32'b10001001000110111100110010110100;
		correct = 32'b10000000000010111000110000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110101100000011000101010010;
		b = 32'b00111001010100110100110011000011;
		correct = 32'b00111000000100000000000001000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000001000100100011100100101;
		b = 32'b10100010111100001100001010011000;
		correct = 32'b10100000001000000100001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111000010101110011000011001;
		b = 32'b01011100011011001111111110011000;
		correct = 32'b00010100000010001110011000011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000100001110010011010110101;
		b = 32'b00010110101101001010010001001000;
		correct = 32'b00000000100001000010010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110110010011000110000011010;
		b = 32'b10011001010100000010000111011101;
		correct = 32'b10000000010000000000000000011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111101101111111101001001100;
		b = 32'b11000000111000011000101001111011;
		correct = 32'b00000000101000011000101001001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100111110100001110101100100;
		b = 32'b10101011011101000011110111111001;
		correct = 32'b00100000011100000001110101100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101000000001101101110101011;
		b = 32'b00001101101101101011110110110111;
		correct = 32'b00000101000000001001100110100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111110100101010110010000101;
		b = 32'b10110110100111001010010110101101;
		correct = 32'b10110110100100001010010010000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100100010011110101111100101;
		b = 32'b10000100010101101101001000011000;
		correct = 32'b00000100000000001100001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011011001000100100000000101;
		b = 32'b00101101101111110100011110000000;
		correct = 32'b00101001001001000100000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001110010111011000110000110;
		b = 32'b11000100111110111101010100001010;
		correct = 32'b01000000110010111001000100000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011101010001100110010000011;
		b = 32'b00100110101100011000010000010010;
		correct = 32'b00000010101000001000010000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111001110010010000010111111;
		b = 32'b11101001010000001011101100110010;
		correct = 32'b01000001000000000010000000110010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010110110010010010000111001;
		b = 32'b11000100111000111010111010000101;
		correct = 32'b00000000110000010010010000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101000100101010101110101110;
		b = 32'b01010001100010111110001001000100;
		correct = 32'b01010001000000101010001000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100001010100011011111101000;
		b = 32'b00011101100111000111111111000011;
		correct = 32'b00010100000010000011011111000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001010100011110110000111101;
		b = 32'b01111011000011100001000101100111;
		correct = 32'b01100001000000000000000000100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010011010111001011110111111;
		b = 32'b10001110000000110101010011010101;
		correct = 32'b10001010000000110001010010010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100100110001011110111111111;
		b = 32'b00011010001100011111101001000001;
		correct = 32'b00000000000100001011100001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011111000010011000011101101;
		b = 32'b00111001011111111011111111100010;
		correct = 32'b00111001011000010011000011100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011110101010101100001111011;
		b = 32'b01101111110010000000111000010011;
		correct = 32'b01001011110000000000100000010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011001001011111001000101000;
		b = 32'b01100111011101101110010101111011;
		correct = 32'b01000011001001001110000000101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111000101111010100101001111;
		b = 32'b10000000011100110100101010100100;
		correct = 32'b00000000000100110000100000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111010011100111001000001000111;
		b = 32'b01010010100000101011000100000010;
		correct = 32'b01010010000000101001000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001111010101101100100000101;
		b = 32'b01010100101011101011101100010001;
		correct = 32'b00000000101010101001100100000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000111100101011111001010110;
		b = 32'b11000111010001100100000110010001;
		correct = 32'b00000000010000100000000000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010001001111101110011110000;
		b = 32'b11110001100101100111111111000010;
		correct = 32'b01110000000001100101110011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101110000010110000110111100;
		b = 32'b10001110000100011010001101011010;
		correct = 32'b00001100000000010010000100011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101001111100101000000010000;
		b = 32'b11110101010011111101111101001111;
		correct = 32'b00110101000011100101000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110000111011000001000111010;
		b = 32'b01000110110101001010011110100111;
		correct = 32'b00000110000101001000001000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111001101001110000000010110;
		b = 32'b00001001000110110010111110011011;
		correct = 32'b00000001000100000010000000010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101011000110100011000100000;
		b = 32'b01001001111001010111000001100100;
		correct = 32'b01000001011000010100000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100110100011101110101111110;
		b = 32'b00001111110001100100101010011000;
		correct = 32'b00000100110000000100100000011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010011000111101010101010011;
		b = 32'b11010001001111100101110100110110;
		correct = 32'b10000000001000100101010100010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110101110010101100100110110;
		b = 32'b10000110001001100011001101111000;
		correct = 32'b00000110001000000001000100110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010011000011011101001000101;
		b = 32'b01000001101110100110000101110011;
		correct = 32'b00000000001000000010000001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100101100010101000100000111;
		b = 32'b11011100000011001111100010000001;
		correct = 32'b11001100000000000101000000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000000001100000000000001100;
		b = 32'b00001111111101011100110111011101;
		correct = 32'b00000000000001000000000000001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001101011011011010111010111;
		b = 32'b11010111100101110001000110101100;
		correct = 32'b00000001100001010001000110000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011011100011000011000101110;
		b = 32'b10100000010000001000010000000010;
		correct = 32'b00100000010000001000010000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101111110101010010000110111;
		b = 32'b10111010011110000110111011001111;
		correct = 32'b10100000011110000010010000000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111111100001001000001101110;
		b = 32'b10000110001001000001010010111101;
		correct = 32'b10000110001000000001000000101100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010000011001011110111010110;
		b = 32'b11000101001001011000001111001101;
		correct = 32'b01000000000001001000000111000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110110010001111010100100010010;
		b = 32'b10110100001111011111100100000100;
		correct = 32'b00110100000001011010100100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000000000001011100100110101;
		b = 32'b00011110011000001000001000100011;
		correct = 32'b00011000000000001000000000100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101010011000000001110101101;
		b = 32'b10010011010000100000110011001011;
		correct = 32'b00010001010000000000000010001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000101110100101001111101101;
		b = 32'b00111111110110110100011101111111;
		correct = 32'b00101000100110100100001101101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100111010010000001011001110;
		b = 32'b10111111100101000111000100110000;
		correct = 32'b10011100100000000000000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111000111011100001100001100;
		b = 32'b01100110111011100001110010001001;
		correct = 32'b01100110000011000000000000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011100100010101100100010101;
		b = 32'b11110101101100001100001000010010;
		correct = 32'b01100001100100000100000000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001111011001110011001011011;
		b = 32'b01011110001010001111111100000111;
		correct = 32'b00001000001010001110011000000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101100110011010101101110111;
		b = 32'b01011100010000010011111111100010;
		correct = 32'b01010100000000010010101101100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110110001001100010001001001;
		b = 32'b00101101001111110110001110010110;
		correct = 32'b00101100000001000100000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000111100000110000001110100;
		b = 32'b10011000001001000001100010011111;
		correct = 32'b10010000001000000000000000010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001111110001101001000011111;
		b = 32'b01000101010100110010111100110001;
		correct = 32'b01000001010100000000001000010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111011100010110001110011111;
		b = 32'b01110100110111011110101011000110;
		correct = 32'b00110100010100010110001010000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000000001011001011010110010;
		b = 32'b11011100001001110011010111000101;
		correct = 32'b00010000000001010001010010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110100100001100110010011011;
		b = 32'b11000000000110011010111110010111;
		correct = 32'b10000000000100001000110010010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111010111011110111010010011;
		b = 32'b01010000011011010111101000110011;
		correct = 32'b01000000010011010110101000010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011011011111100010001110001;
		b = 32'b01000010000001101101100100010011;
		correct = 32'b01000010000001101100000000010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100001011110011010110010010;
		b = 32'b01101111110000100100001010110001;
		correct = 32'b00000100000000100000000010010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111100101101011100101001101;
		b = 32'b10100110011010111010100101100001;
		correct = 32'b00000110000000101010100101000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000110110011010011000011100;
		b = 32'b01011111010001000110111100110101;
		correct = 32'b00001000010000000010011000010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011101001011100010000110101;
		b = 32'b10001100001001011001110010110101;
		correct = 32'b00001000001001011000010000110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111011100101111100101101101;
		b = 32'b01100111110000001100011110100000;
		correct = 32'b00000111010000001100000100100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010011100001000010000001101;
		b = 32'b01111101111101101100001000110010;
		correct = 32'b00010000011100001000000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001101011101101000010010001;
		b = 32'b01000111011001011010110000110101;
		correct = 32'b00000001001001001000000000010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100110111011100010000100000;
		b = 32'b11110101001011101011001001100001;
		correct = 32'b01000100000011001000000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001111110000101110111011111;
		b = 32'b00111011001101100111111111100010;
		correct = 32'b00110001001100000101110111000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101110011100000011100101010;
		b = 32'b10100010000011100100101001001001;
		correct = 32'b10000000000011100000001000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001111000111100111111110000;
		b = 32'b00011010011101011101011010001111;
		correct = 32'b00000000011000011100011010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100011111110011111111101000;
		b = 32'b01100100000000011101011001111100;
		correct = 32'b01000100000000010001011001101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100101100010010001001010111;
		b = 32'b10001010001110101110010001110010;
		correct = 32'b10000000001100000010000001010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111011100100000001110110000;
		b = 32'b10010111010000111010100101010011;
		correct = 32'b10010111010000100000000100010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000010100101011000001101010;
		b = 32'b11000000010110101100001000100101;
		correct = 32'b01000000010100101000000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000000101111111001000101011;
		b = 32'b00001111001001100011000100000111;
		correct = 32'b00000000000001100011000000000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111001001000100110001111111;
		b = 32'b10001100010100110110101111111101;
		correct = 32'b00000100000000000100100001111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000110010010000000110110100100;
		b = 32'b01010110000001110101101111100111;
		correct = 32'b00000110000000000000100110100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111010111010000110110110010;
		b = 32'b00001110001001110000111101001011;
		correct = 32'b00001110000001010000110100000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101101100110101100111001010;
		b = 32'b10010110110010100010001111100101;
		correct = 32'b10010100100000100000000111000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001101101000000010101110101;
		b = 32'b01111110010110110000010110100101;
		correct = 32'b01101000000100000000010100100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000010010101110011010110110;
		b = 32'b11010001110010101010100110010111;
		correct = 32'b01000000010010101010000010010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011101001101101100000101000;
		b = 32'b00001011000001101011000110010100;
		correct = 32'b00001011000001101001000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110000011110001100000011011;
		b = 32'b10110001110011011101111101110010;
		correct = 32'b10010000000011010001100000010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100110010011010011110010110;
		b = 32'b01001011000010001010110011110110;
		correct = 32'b00001000000010001010010010010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011111001111001110011001000;
		b = 32'b00110000110000111011011101000011;
		correct = 32'b00000000110000111001010001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001011011100101000010000111;
		b = 32'b10110101100010001111100111100101;
		correct = 32'b10000001000010000101000010000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010001111001000111000100110;
		b = 32'b11110011000011010110101101110000;
		correct = 32'b10110010000011000000101000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100110111101110101010101100;
		b = 32'b10011100110110010110100010011010;
		correct = 32'b10001100110110000110100010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111010100011111010110111110;
		b = 32'b01000011111111000100110111101110;
		correct = 32'b00000011010100000100010110101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110001111101011010011000110;
		b = 32'b01101011000011110100101000110011;
		correct = 32'b00100010000011100000000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110101111101001110101001000;
		b = 32'b01100101000100000011110000101110;
		correct = 32'b00100100000100000001110000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101011000011001010100000111;
		b = 32'b01010110101011100011111100100001;
		correct = 32'b00010100001000000001010100000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001101101011111010110010100;
		b = 32'b10001111011010100000100101000100;
		correct = 32'b00001001001000000000000100000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101101010100110110101010110;
		b = 32'b00110100000101001000100000010000;
		correct = 32'b00110100000000000000100000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110100010001101011000011100;
		b = 32'b01010001011011101001001110010010;
		correct = 32'b01000000000010001001001000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110001001101010101110011101;
		b = 32'b00011011011000110001111110000111;
		correct = 32'b00000010001000100000101110000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111110001010111001011000001;
		b = 32'b10000101100000100011111100001110;
		correct = 32'b10000101100000000011001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100011111111111000111010000;
		b = 32'b11001000010101000000100110000011;
		correct = 32'b10001000010101000000000110000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101001100011000101110111010;
		b = 32'b11111001111100001000101010001100;
		correct = 32'b01110001001100001000101010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110000011100001000111011011;
		b = 32'b00001000001111000110110101000000;
		correct = 32'b00000000000011000000000101000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010010111101101010111110111;
		b = 32'b00011111101011001010100001000000;
		correct = 32'b00001010000011001000000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011011101000111001101101101;
		b = 32'b00111010000111010101101101111100;
		correct = 32'b00100010000101000101001101101100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010110111100011100110010011;
		b = 32'b00000111100111110000100101010000;
		correct = 32'b00000010100111100000100100010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101001010101101100100011010;
		b = 32'b01010111010000100101110100110001;
		correct = 32'b01010101000000100101100100010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101001101101011010101101111;
		b = 32'b00001011111110000010101101010110;
		correct = 32'b00001001001100000010000101000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100010000000000010110111100;
		b = 32'b10010010011000100100111011010111;
		correct = 32'b00010000010000000000010010010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101011110001111100101011101;
		b = 32'b01001111001010000110100111010011;
		correct = 32'b00000101001010000110100101010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110000010101111101011011110;
		b = 32'b01010111101001111111011100110010;
		correct = 32'b01010110000000101111001000010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101010110111001010110001110;
		b = 32'b00010011001010011011001010101001;
		correct = 32'b00000001000010011001000010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011010110001101001001111010;
		b = 32'b00110100110001110010011001010101;
		correct = 32'b00000000010000000000001001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011100011110000011011001111;
		b = 32'b11001110101010110000111011110001;
		correct = 32'b01001010100010110000011011000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001001000101111000101011101;
		b = 32'b10101111110000001110001010000001;
		correct = 32'b00000001000000001110000000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100101011101101101010110000;
		b = 32'b11100001010111110011010101111000;
		correct = 32'b10100000000011100001000000110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111010000011110011100100101110;
		b = 32'b01000010001111110000011110010000;
		correct = 32'b01000010000011110000000100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011111111110000111110010011;
		b = 32'b01110110100111000110010000101001;
		correct = 32'b01100010100111000000010000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100110000100011011110101000;
		b = 32'b10110111101000001100010011111101;
		correct = 32'b10010100100000000000010010101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111100111110011101100101011;
		b = 32'b00000111100001110011100010011100;
		correct = 32'b00000111100001110011100000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001011011000001001001001001;
		b = 32'b10001000101111001000010011000100;
		correct = 32'b10001000001011000000000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010101111111101001110100101;
		b = 32'b10111011110010100101111001010100;
		correct = 32'b10101010100010100101001000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110100101001011110001100111;
		b = 32'b00010000100110100111101110110101;
		correct = 32'b00010000100100000011100000100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111110101110100010001000100;
		b = 32'b00111011011010110011010011100010;
		correct = 32'b00110011010000110000010001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001101001010011111100010001;
		b = 32'b10010110010111011111001111111010;
		correct = 32'b00000000000001010011001100010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001111010011111111100101011;
		b = 32'b11111000110110101001001011101110;
		correct = 32'b00010000110010001001001000101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101011100011001110000001000;
		b = 32'b11100111001001111000110111000100;
		correct = 32'b10000101001000011000110000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011001011001110000111001011;
		b = 32'b01000001101100110101110111000000;
		correct = 32'b01000001001000000100000111000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101011100010100011101010111;
		b = 32'b01001011100111010000011110011010;
		correct = 32'b00001001000100010000011100010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001000000000010001111111110;
		b = 32'b11111010010110010110011011001110;
		correct = 32'b11101000000000000010001011001110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111110100110100111000001110;
		b = 32'b11101010111001111110011111001001;
		correct = 32'b01101010110000110100011000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011110011100001010010010000;
		b = 32'b01101101011100111001110111001101;
		correct = 32'b00001001010000100001010010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011100000100100101101100101;
		b = 32'b00100010100010011000000000011001;
		correct = 32'b00000010100000000000000000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111101011011111011011000111;
		b = 32'b11000110000100110001100001100011;
		correct = 32'b10000110000000010001000001000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111001101110011000000100000;
		b = 32'b00111101010110101111101010001011;
		correct = 32'b00111101000100100011000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100001010001110011110100001;
		b = 32'b01100010010011001101111100100010;
		correct = 32'b01100000000010001100011100100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010110001010110000001011001;
		b = 32'b11100000111101000010111011010101;
		correct = 32'b11000000110001000010000001010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010001111000010100000100010;
		b = 32'b11100000111010010100101011000100;
		correct = 32'b11100000001010000000100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100101000100001111011010001;
		b = 32'b11011110001110100001000001101101;
		correct = 32'b01011100001000100001000001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101011101001010010110010011;
		b = 32'b01100011111110000011110010000100;
		correct = 32'b00000001011100000010010010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110011001111100011110110110;
		b = 32'b01001010100110010111010011011001;
		correct = 32'b00001010000000010100010010010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110111111100000011111000010;
		b = 32'b11101011011000101100110010000110;
		correct = 32'b10001010011000100000010010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110101001010100011101100100;
		b = 32'b00101111101100001001010000110001;
		correct = 32'b00100110101000000000010000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111000111000110011111111100;
		b = 32'b01000110110000100001110011010111;
		correct = 32'b01000110000000000000010011010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000100101011100001000000010;
		b = 32'b11110110110010100001010000010101;
		correct = 32'b11010000100000000000000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000100100011101000001110111;
		b = 32'b11011011111000001011010100101110;
		correct = 32'b11010000100000001001000000100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001110001110110111011000101;
		b = 32'b10001010010011101111100010101101;
		correct = 32'b00000000010001100110100010000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111010110000111100001000100;
		b = 32'b01101001010111100010001101101011;
		correct = 32'b00000001010110000010000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111110010101110110000010100;
		b = 32'b11111110110110111000001101100101;
		correct = 32'b10100110110010101000000000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001001101011001011100000000;
		b = 32'b11011010001001010000101111111110;
		correct = 32'b11000000001001010000001100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101110000001000110110000110;
		b = 32'b11110001100000000010010010010000;
		correct = 32'b01010001100000000000010010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111100010011111010010000000;
		b = 32'b10111100001101111100110011000110;
		correct = 32'b10100100000000011100010010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100000001000100000000100101;
		b = 32'b10000001000011000010100111101001;
		correct = 32'b00000000000001000000000000100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110101111001001000011101000;
		b = 32'b10000100100110110111001100110010;
		correct = 32'b10000100100110000001000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010101011011001011000000101;
		b = 32'b10110010111110110111011001110110;
		correct = 32'b10110010101010010001011000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000001000001101110010010001;
		b = 32'b10100110110011111010011100100100;
		correct = 32'b00000000000000001000010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010011100011000111100110100;
		b = 32'b10011001000100111110101111000100;
		correct = 32'b10010000000100011000101100000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110001110010101111110110000;
		b = 32'b11101010000100001101110110101111;
		correct = 32'b01101010000100000101110110100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011011011001001100001111001;
		b = 32'b10110011001000101011000000010001;
		correct = 32'b00110011001000001001000000010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111000000000100100111101001;
		b = 32'b10111000101000111111001111101011;
		correct = 32'b10101000000000000100000111101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011000100001001110011010101;
		b = 32'b11111011010111101001110011001000;
		correct = 32'b11111011000100001001110011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101100001001010011110011001;
		b = 32'b11000101100110011001001110011101;
		correct = 32'b00000101100000001000001110011001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010001100001010100100010010;
		b = 32'b00111010111100010100111010110110;
		correct = 32'b00000010001100000000100000010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101110101011001011001010001;
		b = 32'b11011011111101000010011101110011;
		correct = 32'b10001001110101000000011001010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101000101110110110101011110;
		b = 32'b01110011111111100011111101011010;
		correct = 32'b01110001000101100010110101011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010000110100101010101010101;
		b = 32'b10101010000010110000001011111000;
		correct = 32'b10101010000010100000000001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010010100000001111001010111;
		b = 32'b11011101001001010011111110110010;
		correct = 32'b00000000000000000001111000010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010011100001100111101101111;
		b = 32'b01111101111111010001011011001000;
		correct = 32'b01001000011100000000011001001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011001100011000110100100000;
		b = 32'b11011110101010000100100100010100;
		correct = 32'b01000010001000000000100100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101001110110011000110011000;
		b = 32'b01110010111101010110000001111001;
		correct = 32'b00110000001100010010000000011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111010000110111100000100110;
		b = 32'b11010111100000111011001101000101;
		correct = 32'b11010111000000110011000000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010010000001001111111011100;
		b = 32'b11111000101001010100010000101110;
		correct = 32'b01011000000000000000010000001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101010001000000101011000010;
		b = 32'b10101100001111010100000110001011;
		correct = 32'b10101100000001000000000010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011001000100010010011110010;
		b = 32'b11101011011110111000110010001110;
		correct = 32'b01000011001000100000010010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101000100100110010001011011;
		b = 32'b11101001110000010011010000000011;
		correct = 32'b01000001000000000010010000000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001101100100000101000001011111;
		b = 32'b01101010111001111011010111111010;
		correct = 32'b00001000100000000001000001011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000100111101110000110010111;
		b = 32'b11001000100001010110110101101000;
		correct = 32'b10000000100001000110000100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011110101101001000100101001;
		b = 32'b10000100000010001001010100100110;
		correct = 32'b00000000000000001001000100100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111000001111110011100101111001;
		b = 32'b01100100010111100110100110000001;
		correct = 32'b01100000000111100010100100000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100000101100110101101110000;
		b = 32'b01111000001011000010111100001110;
		correct = 32'b00111000000001000010101100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000100010000100000010000000;
		b = 32'b01011001000100010011001111011110;
		correct = 32'b01011000000000000000000010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000101100011111111000111011;
		b = 32'b01010111111011100001111111100000;
		correct = 32'b01000000101000000001111000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011110101101001011000001000;
		b = 32'b01111110101111110101001111111111;
		correct = 32'b00100010100101100001001000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100100101111110000101000000;
		b = 32'b00010010001101011001101011010110;
		correct = 32'b00000000000101011000000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001110101011111011001110010;
		b = 32'b00101001110001100011100010000010;
		correct = 32'b00100001110001000011000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011111010111010000011011000;
		b = 32'b01011001111100011000001000010110;
		correct = 32'b01010001111000011000000000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111010110111000000110100001;
		b = 32'b01111001101011010010011111001101;
		correct = 32'b01001001000010010000000110000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110111001111110010110000111;
		b = 32'b11011101111001100100000001110011;
		correct = 32'b01010100111001100100000000000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101110001011010111101010100;
		b = 32'b10011010110101111110100010100010;
		correct = 32'b00000000110001011010100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111111110111001011000110111;
		b = 32'b00100010000010000001100010110111;
		correct = 32'b00000010000010000001000000110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100011001111110110101010110;
		b = 32'b00000101011111011100001110000110;
		correct = 32'b00000100011001011100000100000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111110110111101110100111001;
		b = 32'b11011100000100101001101010101011;
		correct = 32'b01011100000100101001100000101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001100110101001000001010111;
		b = 32'b11011110000100000101110110001010;
		correct = 32'b00010000000100000001000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100101011111000110000011111;
		b = 32'b11001111110101011101011101110011;
		correct = 32'b11001100100001011000010000010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110010110011001011111111111;
		b = 32'b00101010000110100110000110001111;
		correct = 32'b00100010000110000000000110001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001101001111111111111000100;
		b = 32'b01101001001100000011000011110101;
		correct = 32'b01100001001000000011000011000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101111111001101011101111001;
		b = 32'b10000010000111000011110111100111;
		correct = 32'b00000000000111000001010101100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111111111011011100000100001;
		b = 32'b00100011111101101111000010011000;
		correct = 32'b00100011111101001011000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011111000111101100110100011;
		b = 32'b10010010000100001101000010100110;
		correct = 32'b00000010000000001101000010100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000010000101000100110011001110;
		b = 32'b01011010111010101011101010011001;
		correct = 32'b00000010000000000000100010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011100000010000011011000101;
		b = 32'b00011001000111011101010111010110;
		correct = 32'b00001001000000010000010011000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110011101101000011111001101;
		b = 32'b11011010110010010011100101101011;
		correct = 32'b10011010010000000000000101001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011111001100001101001011010;
		b = 32'b00100111011011111100001000001101;
		correct = 32'b00000011011001100000001000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001001111110101101000000000;
		b = 32'b01010111101011110111111010111110;
		correct = 32'b01010001001011110101101000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011001001011001110110111000;
		b = 32'b00111111110101101110001011100100;
		correct = 32'b00100011000001001000000010100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101101100000100001110011110;
		b = 32'b00101111111010101111111000110010;
		correct = 32'b00100101101000000100001000010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101011110010000000000001100;
		b = 32'b11101101000001100100011111111110;
		correct = 32'b11000101000000000000000000001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011110111001000010111100011;
		b = 32'b01111011010011110110000111101001;
		correct = 32'b00101011010011000000000111100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000111001101001101011011101010;
		b = 32'b00111110101100001110000010000011;
		correct = 32'b00000110001100001100000010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001110010101011001011001011;
		b = 32'b00110111010101010101100010011001;
		correct = 32'b00110001010000000001000010001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000000001110011101000011000;
		b = 32'b11011101100010111011110011000110;
		correct = 32'b01010000000000110011100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111011100010110011101100110;
		b = 32'b00000111110000110111000111010110;
		correct = 32'b00000111010000010110000101000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100011010100111110010101111;
		b = 32'b01101010100000000110110010011011;
		correct = 32'b00000000000000000110110010001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001101110001101001111111101;
		b = 32'b10111001101000100000101110001100;
		correct = 32'b10111001101000000000001110001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100010111100001001001010111;
		b = 32'b11101011001011000010000000001101;
		correct = 32'b00100000000011000000000000000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100111110010101100001010011;
		b = 32'b11001000101100000101001100111111;
		correct = 32'b10001000101100000101000000010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100101110101101111100000111;
		b = 32'b10100110110110011100011110101101;
		correct = 32'b10000100100110001100011100000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101010111101111100000010100;
		b = 32'b00010111110011011110110101110011;
		correct = 32'b00010101010011001110100000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000110000101100010111100010;
		b = 32'b00101100100010010111110101001000;
		correct = 32'b00100000100000000100010101000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100101000100011000101010101;
		b = 32'b11101001001110111001111000100011;
		correct = 32'b00101000001000100001000000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011001001100100001111100100;
		b = 32'b00011100001111111111000000001110;
		correct = 32'b00000000001001100100000000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110010111011011100001000001;
		b = 32'b01110000001101100101000001000010;
		correct = 32'b00110000000101000001000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010101110101100001101101001;
		b = 32'b01010111100100111100110110001100;
		correct = 32'b01010010100100101100000100001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101110000110101100101101111;
		b = 32'b10101100111000000110000100011100;
		correct = 32'b10100100110000000100000100001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001101010010100111000100010;
		b = 32'b01111010011011101101110010110100;
		correct = 32'b01011000001010000100110000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010001011010001110110101010;
		b = 32'b10111100010111101011010111000010;
		correct = 32'b10000000000011000001010110000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011000100010111111100011101;
		b = 32'b10110000001000011101010101111010;
		correct = 32'b00110000000000010101010100011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000011011111100010100111100;
		b = 32'b11101010001011001001110100010010;
		correct = 32'b01001000001011001000010100010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010110010010110010001011001;
		b = 32'b11101001110000000111110010101000;
		correct = 32'b01101000110000000110010000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110010011000000001000000110;
		b = 32'b11100111110110011010000010101010;
		correct = 32'b00000110010010000000000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010011101000110101011101110;
		b = 32'b01000000111000110000101110001100;
		correct = 32'b00000000011000000000101010001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110110001110101100100101101;
		b = 32'b11100011111110101010101011011100;
		correct = 32'b11000010110000100000100000001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110111011010111000110100110;
		b = 32'b10101111101001101100010111100010;
		correct = 32'b10100110101001000100000110100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010101111100011010011100010;
		b = 32'b01011011000101010101001100100011;
		correct = 32'b01000010000101000001000000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100011010010111101110000110;
		b = 32'b01100110111111110001001001011011;
		correct = 32'b00100100011010010001001000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111110011001011010101101110;
		b = 32'b01111010101001000000100010010011;
		correct = 32'b00010010100001000000000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101110100100101000010010111;
		b = 32'b10011100101000100000101100110111;
		correct = 32'b00001100100000100000000000010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110111011011010110011000100;
		b = 32'b01100010111100011110110010101011;
		correct = 32'b00000010111000011010110010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011111001100101010010000001;
		b = 32'b00001110100110000010000110100010;
		correct = 32'b00001010100000000000000010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111011000001100111010001011;
		b = 32'b01110011011110001100000001001000;
		correct = 32'b01100011011000001100000000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111111010110100100110000110;
		b = 32'b01001001000000001001101001100100;
		correct = 32'b01001001000000000000100000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001100101110010100101000101;
		b = 32'b11011001110110001110011110011000;
		correct = 32'b00010001100100000010000100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010111011010001011011101101;
		b = 32'b01011000101101101101001001101101;
		correct = 32'b01001000101001000001001001101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011110101101111110110000000;
		b = 32'b11111100101010000110110001010100;
		correct = 32'b01001000100000000110110000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001100110101000000101000011;
		b = 32'b00011001101011010111000111111011;
		correct = 32'b00011001100010000000000101000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000101101011111100001001001;
		b = 32'b11101001111100000100111000110000;
		correct = 32'b01000000101100000100100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000101111101001000101101000;
		b = 32'b11011111110011010110010101111100;
		correct = 32'b11000000100011000000000101101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011111001101011110011110111;
		b = 32'b00100010011000011100101111010100;
		correct = 32'b00100010011000001000100011010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101101110011011111010101010;
		b = 32'b11101111100101001010101110101100;
		correct = 32'b10101101100100001010101010101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000100011110100111011010001;
		b = 32'b01111110001000011010001001000011;
		correct = 32'b01010000000000010000001001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011111111101010001010100110;
		b = 32'b11100001010110110000011000010000;
		correct = 32'b00000001010110100000001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011010111110011000101101110;
		b = 32'b10011100101000101111100010101110;
		correct = 32'b10010000000000100011000000101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100111100000011010110101011;
		b = 32'b00100101011100011011110100010100;
		correct = 32'b00000100011100000011010100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101010101110001111110110011;
		b = 32'b00111000001011010111110101111001;
		correct = 32'b00011000000001010001110100110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101111101001011111010000110;
		b = 32'b11001010100011011001010101011100;
		correct = 32'b00000000100001001001010000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001000110000010000000110011;
		b = 32'b01110001000010100000100110110001;
		correct = 32'b01000001000010000000000000110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101010101010000010010001110;
		b = 32'b10111111110100011000011010101010;
		correct = 32'b00110101010100010000010010001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000011110011110010001100111;
		b = 32'b10111001110000001100110011100101;
		correct = 32'b10100000010000001100010001100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001111001001111011110101011;
		b = 32'b10100011001010111001000110010110;
		correct = 32'b00100001001000001001000110000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001101001000000111011001101;
		b = 32'b00100100010011101111100000001110;
		correct = 32'b00100000000001000000100000001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100100101011100101101010001;
		b = 32'b10100111011100011001000001110111;
		correct = 32'b00100100000100011000000001010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000101111101001111001000100;
		b = 32'b01010010010001010111110101111010;
		correct = 32'b00010000000001000001110001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001001000110000110001010100;
		b = 32'b10000001101010011010100110111101;
		correct = 32'b10000001001000010000100000010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111100001101000111000000100;
		b = 32'b10101100010011111011111110010001;
		correct = 32'b10101100000001101000111000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001101110001011100110101011;
		b = 32'b01000110001111100100010101000010;
		correct = 32'b01000000001110000000000100000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110010100010100111100000001;
		b = 32'b01101110001100001111100101111011;
		correct = 32'b01001110000100000100100100000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000011110001010111010011101;
		b = 32'b00000010010011010111101101010110;
		correct = 32'b00000000010010000010101000010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101110000100010110101001000;
		b = 32'b11000100001100101101110101110111;
		correct = 32'b10000100000000100000110101000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101101010100101110011101100;
		b = 32'b00111110011010100100100010110110;
		correct = 32'b00010100001010100100100010100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000011001000110011101010100;
		b = 32'b00110100100111110101111110000001;
		correct = 32'b00100000000001000100011100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101011101110011101000110011;
		b = 32'b00111110011110010100010011100100;
		correct = 32'b00110100011100010000000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100011001010111010111111101;
		b = 32'b00001001010000101101001001000011;
		correct = 32'b00000000010000000101000001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110111110010001111111101111;
		b = 32'b11100110111111001001100111000000;
		correct = 32'b11100110111110000001100111000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011010011100101110010010110;
		b = 32'b00001110000110000000101001110100;
		correct = 32'b00001010000010000000100000010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110000001111100000110101111;
		b = 32'b11100010101001100110010001110000;
		correct = 32'b11100010000001100100000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110011011010011001001100101;
		b = 32'b11110000101110111001010011100100;
		correct = 32'b01100000001010010001000001100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001001011010101001110101101;
		b = 32'b01010010111010100110000011000100;
		correct = 32'b01010000001010000100000010000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011011011101010001001110001;
		b = 32'b00100101100101101100101101101011;
		correct = 32'b00000001000001101000001001100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011011010010111101110000001;
		b = 32'b00100111100110011001011010000110;
		correct = 32'b00100011000010010001001010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010101101010101100100111110;
		b = 32'b01110110110100011001011110111010;
		correct = 32'b01110010100100010001000100111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000111110010001100100001110101;
		b = 32'b00111111000001100000010101000011;
		correct = 32'b00000111000000000000000001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010101100010110111101001101;
		b = 32'b01110000110100001001011010111010;
		correct = 32'b00110000100100000000011000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100011101011100110101101111;
		b = 32'b10010010110011110000011111110011;
		correct = 32'b00010000010001010000010101100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000101011101111110000010100;
		b = 32'b00010110100101111111011011001001;
		correct = 32'b00010000100001101111010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010010011101001011111001000;
		b = 32'b10111111100001010111000110000011;
		correct = 32'b00101010000001000001000110000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100001010001000100101101101;
		b = 32'b10111011110011111111101000010101;
		correct = 32'b10111000000010001000100000000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001100101000011001101011101;
		b = 32'b00111000010000010101100011101111;
		correct = 32'b00100000000000000001000001001101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000100100000111011000111111111;
		b = 32'b01011101100001000011100100001010;
		correct = 32'b00000100100000000011000100001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010101011101110110010110100;
		b = 32'b11001011100011000101101000010010;
		correct = 32'b00000010100011000100100000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101001000000100000111110111;
		b = 32'b11100101110011110000100010001010;
		correct = 32'b01000101000000000000000010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010111101101011101010111111;
		b = 32'b01010111110011010100111110000011;
		correct = 32'b00010010110001000000101010000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010001110011000010001011101;
		b = 32'b00011010100111100011001001010101;
		correct = 32'b00011010000110000000000001010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111010001000001110110110011;
		b = 32'b00101110100000010110011101000100;
		correct = 32'b00001110000000000000010100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111111110010000001110111110;
		b = 32'b11001001101011101001110010100011;
		correct = 32'b00000001101010000000000010100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110000111010110001100010001;
		b = 32'b00111001101000110011100100100100;
		correct = 32'b00011000000000010010000100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010010011111010110100110001;
		b = 32'b11111010011001100001011110010001;
		correct = 32'b00111010010001100000010100010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011010000100000010000110010;
		b = 32'b00110000011101111001000101101100;
		correct = 32'b00110000010000100000000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000100110111110010100000001111;
		b = 32'b10101010100111100000010100001011;
		correct = 32'b10000000100111100000000000001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001111011011101000101011010;
		b = 32'b11110011000101011011100111110001;
		correct = 32'b00000001000001011001000101010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011010011001111101110110110;
		b = 32'b11111000101111110101100011000111;
		correct = 32'b00011000000011000101100010000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100000001001000110110000000;
		b = 32'b11101101101000001100111010111010;
		correct = 32'b01101100000000001000110010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110001010111111000100111101;
		b = 32'b01011011101000111100101011000100;
		correct = 32'b01010010001000111100000000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001110001100110110100110111;
		b = 32'b01110010001111010011110111000110;
		correct = 32'b00010000000001000010110100000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111101001000001101110000001;
		b = 32'b10110011101000011011100110111000;
		correct = 32'b00010011101000000001100110000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000111101010010111101010101;
		b = 32'b11101011010110110011010010000100;
		correct = 32'b00001000010100010010010000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000110010001010110000111111;
		b = 32'b00101110100111010001100101100111;
		correct = 32'b00000000100010000000100000100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001101110111000010001110001;
		b = 32'b11000100100110110010101010011100;
		correct = 32'b00000000100110110000000000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010101100001100010100110001;
		b = 32'b00111101101011010110000001100010;
		correct = 32'b00110000101000000100000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100100011100100111011010000;
		b = 32'b10110100000111011001101010011111;
		correct = 32'b00000100000011000000101010010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111010111000011000011011111;
		b = 32'b01000111111100101000100101000110;
		correct = 32'b01000111010100000000000001000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100110100111001100010001010;
		b = 32'b10101100100100010010111011010001;
		correct = 32'b10101100100100010000100010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101110010000000111001001000;
		b = 32'b00011111001100110101111000001101;
		correct = 32'b00000101000000000000111000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001010100110001101110001111;
		b = 32'b01000011001110110100111001111010;
		correct = 32'b00000001000100110000101000001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010001000011111011101101001;
		b = 32'b11000011000100110110001000110111;
		correct = 32'b10000010000000010110001000100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011010101101010111101010110;
		b = 32'b00110111101110100100000111011010;
		correct = 32'b00000011000100100000000101010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110101001010100000011110001;
		b = 32'b01000000100011110110001110000011;
		correct = 32'b01000000100001010100000010000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011001111001101010010101011;
		b = 32'b01101011010010111110111001001001;
		correct = 32'b01001011000010001100010000001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000101110001111110110110110;
		b = 32'b01010001011001100000001110111000;
		correct = 32'b00000000001000000000000110110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010010010111110100100101011;
		b = 32'b10010010100111101010010110110001;
		correct = 32'b10010010000010101010000100100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101110011100110111101100000;
		b = 32'b00001011001111001000111101100001;
		correct = 32'b00000001000011000000111101100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010000000110011100111010010;
		b = 32'b00000010001110100100101100100011;
		correct = 32'b00000010000000100000100100000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001111111001110100010001001;
		b = 32'b01010010101101001101100101100000;
		correct = 32'b00010000101101001100100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110001100101111001001100101;
		b = 32'b11111010010101011000010001000010;
		correct = 32'b00010010000100001000000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110111001100010101000001011;
		b = 32'b10011110011101111010011101111110;
		correct = 32'b00010110011001100010001000001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011110101001000001100000010;
		b = 32'b00100110100001110011111001101111;
		correct = 32'b00000010100001000000001000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000110011001110001101001010;
		b = 32'b10110101011111010110001101011011;
		correct = 32'b10100000010011000110001101001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110110101111001110011110110;
		b = 32'b10001101001010101001100000010111;
		correct = 32'b10001100000000101001100000010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001010111001011100100101101;
		b = 32'b10110101100110001000000010011010;
		correct = 32'b00110001000110001000000000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101000100001111111100010001;
		b = 32'b01000101000111100100111111011011;
		correct = 32'b01000101000100000100111100010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000010101010110011001010100;
		b = 32'b01101101001110100011001100010011;
		correct = 32'b01001000000100000010001000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011111001011011101000110000;
		b = 32'b00100100110100100111010110100101;
		correct = 32'b00100000110000000011000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010110111101101010110010100;
		b = 32'b01101000000111110101000010110000;
		correct = 32'b00001000000111100101000010010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101000111010100101101000010;
		b = 32'b00000110110110100101000011001000;
		correct = 32'b00000100000110000100000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111100111101111110101011101;
		b = 32'b01100101001110000010001111101101;
		correct = 32'b01100101000110000010000101001101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011011011000101111000100011;
		b = 32'b10010100110101110100101111010011;
		correct = 32'b10010000010001000100101000000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101110110011110011110100011;
		b = 32'b00000101011101101101101000010110;
		correct = 32'b00000101010100001100001000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101100100111000100100011001;
		b = 32'b01001010001101001010010100111111;
		correct = 32'b01000000000100001000000100011001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001111001101001010101000101;
		b = 32'b01001011001011001010111010110101;
		correct = 32'b01000001001001001000010000000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101010010000111010110101001;
		b = 32'b11010110101111100101111100111011;
		correct = 32'b11000100000010000101010100101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110111110100111111000000010;
		b = 32'b11101100001100010100000011100000;
		correct = 32'b01100100001100000100000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111000110111010101010100111;
		b = 32'b01010011101011100100000110101010;
		correct = 32'b01000011000010100000000010100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100111011101001010000000100;
		b = 32'b10001011100100010000011101100000;
		correct = 32'b00001000100000000000010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001010001010110111111001110;
		b = 32'b10001000110110100111100001110100;
		correct = 32'b00000000010000000110100001000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011010010000000101101001110;
		b = 32'b00001100001001111001110000011110;
		correct = 32'b00000000000000000000100000001110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110010111100000111011000100;
		b = 32'b01110001011101010100010000110100;
		correct = 32'b00000000010101000000010000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001000011010001010000101111;
		b = 32'b00110011011010100110010100101011;
		correct = 32'b00000001000010000000010000101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001010100000111100111100010;
		b = 32'b10100101010101011010001000111101;
		correct = 32'b00100001010100000010000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000000011000011110100011001;
		b = 32'b11111000100011100011100010111010;
		correct = 32'b11000000000011000011100000011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110010000000000000101001100;
		b = 32'b10011110111100110101110100001111;
		correct = 32'b00011110010000000000000100001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111011000111010100101100101;
		b = 32'b10001010010101010010110111101010;
		correct = 32'b10001010010000010010100101100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100111011100011111001100101;
		b = 32'b10000111011111011000110111100110;
		correct = 32'b00000100011011000000110001100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111001100010001001011001011;
		b = 32'b00000110001001111110110100101111;
		correct = 32'b00000110001000010000000000001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011010111000101001111111110;
		b = 32'b11100011000110011110100000100101;
		correct = 32'b00000011000110000100000000100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100001111101011000100010000;
		b = 32'b01101001001100111000111110011101;
		correct = 32'b01101000001100101000000100010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100001110001011101101000010;
		b = 32'b01110100001110110000111001100111;
		correct = 32'b00010100001110000000101001000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101110001111001101100000101;
		b = 32'b01001111110111000001010001001011;
		correct = 32'b01000101110001000001000000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111101010101110111010100001;
		b = 32'b00000001101000101110000011010101;
		correct = 32'b00000001101000101110000010000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000010000010111111011100010;
		b = 32'b00110110101001011010100001010110;
		correct = 32'b00000000000000010010100001000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001010001101000111010010101;
		b = 32'b01110010011001101100011100000010;
		correct = 32'b00000000010001101000011000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000000100001001000111001100;
		b = 32'b11000011100001100011100011001110;
		correct = 32'b00000000000000000001000011001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010100100101100001000101111;
		b = 32'b10010011101011110101100100011111;
		correct = 32'b10010010100000100100000000001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111000000110010111111101111;
		b = 32'b10100001111100101000010001010100;
		correct = 32'b00000001000000100000010001000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101101100000011111001110101;
		b = 32'b01001001011110111001010000010100;
		correct = 32'b01000001001100000001010000010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100000100010110100110111001;
		b = 32'b01110100101011110000001000101011;
		correct = 32'b00000100000000010000000000101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110110010111001000110111011;
		b = 32'b10111101001110000000100011110110;
		correct = 32'b00111100000010000000000010110010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001011010111011000001101100;
		b = 32'b10110010000000111111111010100010;
		correct = 32'b00000000000000111011000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100110001111101001000011100;
		b = 32'b11100010101010001111011100100001;
		correct = 32'b01000000100000001101001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100010000000101001010101001;
		b = 32'b00111010101111010011011001101101;
		correct = 32'b00101000000000000001001000101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011001010001111010000001110;
		b = 32'b00101101011101010100101010000000;
		correct = 32'b00000001001000000100000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000111011110111011100111001;
		b = 32'b10000101100001100011110001101010;
		correct = 32'b00000000100001100011010000101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011111011001100000010001010;
		b = 32'b01111100110000110000101101011111;
		correct = 32'b00110000110000000000000000001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000010101011001100001000001;
		b = 32'b11101110011110010111100011101110;
		correct = 32'b10000000010100010001100001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110000001110001011111001001;
		b = 32'b10001110110100111100001011000101;
		correct = 32'b00000110000000110000001011000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111100010111110100010110110;
		b = 32'b11111000001001100111001001110001;
		correct = 32'b01100000000000100110000000110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101100001010010000101100011;
		b = 32'b10100100111011111100110100000100;
		correct = 32'b00000100100001010000000100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100001010110101110100010101;
		b = 32'b11001010101100000000100101101100;
		correct = 32'b11000000001000000000100100000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100101101110100100011000001;
		b = 32'b11111100110001101000000111110011;
		correct = 32'b01000100100001100000000011000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101010000100001001100001100;
		b = 32'b01010001100111111111110110111010;
		correct = 32'b01010001000000100001000100001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111000111000000010000111011101;
		b = 32'b00111011111110101100001100101010;
		correct = 32'b00111000111000000000000100001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001101101110010100010110100;
		b = 32'b11010110111101000000001010001010;
		correct = 32'b00000000101101000000000010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110011110110000011011100100;
		b = 32'b10010000110000011010001101000011;
		correct = 32'b00010000010000010000001001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101110100000011111101010011;
		b = 32'b10100011111110011101110010100001;
		correct = 32'b00100001110100000001110000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001101011111100101101011001;
		b = 32'b01110110000111110111010010100110;
		correct = 32'b00100000000011110100000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001111001111010000001110011;
		b = 32'b10010000000011101011000010101001;
		correct = 32'b10010000000001101010000000100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000101010000111000010010000;
		b = 32'b00000000101111011110010001110000;
		correct = 32'b00000000101010000110000000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001111000101000000110011100;
		b = 32'b10000101011000100010001100111101;
		correct = 32'b10000001011000100000000100011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110111110110011111011110110;
		b = 32'b00000010011111000101000111101100;
		correct = 32'b00000010011110000001000011100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100011110111111111001101101;
		b = 32'b01001010110010011010000000100011;
		correct = 32'b01000000010010011010000000100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110011001110000101010011001;
		b = 32'b00111111000000100001110111100000;
		correct = 32'b00001110000000100000100010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111010011100110001010110111;
		b = 32'b11111110110110000001000100001011;
		correct = 32'b11011110010010000000000000000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110011110011110101111010100;
		b = 32'b11001011000011011000111111110010;
		correct = 32'b10001010000010011000101111010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110110100011000001001000000;
		b = 32'b10111100010000110011100101110000;
		correct = 32'b10101100010000010000000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111000011110000001011110011111;
		b = 32'b10110001100011111111111000100011;
		correct = 32'b10110000000010000001011000000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001011010011011010010111111;
		b = 32'b11100000100000110101111101100010;
		correct = 32'b00100000000000010001010000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011011010100100010011001000;
		b = 32'b00100011100010001110100000011000;
		correct = 32'b00100011000010000100000000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011101111101011000111010011;
		b = 32'b01001010001111101010000111011101;
		correct = 32'b00000010001111101010000111010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000011001101110100011111010;
		b = 32'b00101100000101110011101011110110;
		correct = 32'b00001000000001100010100011110010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111010110010111001101111010;
		b = 32'b00100000001100110111111000000101;
		correct = 32'b00100000000100010111001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101101100011110001001011101;
		b = 32'b10110111111100101010010110001010;
		correct = 32'b10100101101100001010000000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110110011111000101101100101;
		b = 32'b11110111100001100010101110110111;
		correct = 32'b10100110100001100000101100100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110110111000011010011001011;
		b = 32'b01000101100111011101100010101100;
		correct = 32'b00000100100111000001000010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001011101101100100100101111;
		b = 32'b01111000100000100000101101111011;
		correct = 32'b00000000000000100000100100101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111010101000110000010111011;
		b = 32'b11100101011001110101100000011010;
		correct = 32'b01000101010001000100000000011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100101010001010100101010010;
		b = 32'b11100000010100111000100011110010;
		correct = 32'b00000000000000001000100001010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001011110010011111100011111;
		b = 32'b00111110101001111101011111001001;
		correct = 32'b00010000001000010001011100001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011010101100101110000010010;
		b = 32'b11000000100010011101011010101111;
		correct = 32'b10000000000000000101010000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010001001000100111110101000;
		b = 32'b01001001001101111011110110110001;
		correct = 32'b01001000001001000000110110100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111000011100110111010101010010;
		b = 32'b10110101010111010101110111011111;
		correct = 32'b10110000010100010101010101010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110000010111110101001001101;
		b = 32'b11101011010011001001001000101110;
		correct = 32'b10101010000010001000001000001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110110001101111111001010100;
		b = 32'b01000101111111000111010110010111;
		correct = 32'b01000100110001000111010000010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011100001101011111110110110;
		b = 32'b11111001001010111101010011101010;
		correct = 32'b00111001000000101001010010100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110000000111101101111010010;
		b = 32'b10001110000000010000111000000110;
		correct = 32'b10001110000000010000101000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001110101110001100001000011;
		b = 32'b11000101000111101110111110010000;
		correct = 32'b11000001000101100000100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010010110110001000000000110;
		b = 32'b10011110000110100111100001100010;
		correct = 32'b00000010000110100001000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110111111011001010000001010;
		b = 32'b10001110001000110001000111000110;
		correct = 32'b10001110001000010001000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011101000000010001010011000;
		b = 32'b01001000110001011111110111100110;
		correct = 32'b01000000100000000010000010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111010011111101011010100111;
		b = 32'b01100001110101011001101111000110;
		correct = 32'b00000001010001011001001010000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100000101101111111010000111;
		b = 32'b00101010110101000101000111110101;
		correct = 32'b00001000000101000101000010000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111010010000000010110110000;
		b = 32'b00011110001001100000010101011100;
		correct = 32'b00011110000000000000010100010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101110001001010010000101100;
		b = 32'b11111110101000101001111111100001;
		correct = 32'b01111100100000001000010000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011111101101110011011101001;
		b = 32'b00101000011011001010100101000111;
		correct = 32'b00100000011001001010000001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000001101110101011001001000;
		b = 32'b01000110001101100111100111010000;
		correct = 32'b00000000001101100101000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001000110100111010001110011;
		b = 32'b00011110011001011100111111111101;
		correct = 32'b00011000000000000100010001110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110100010011000001110100000;
		b = 32'b10001000011111101100110111110111;
		correct = 32'b10000000000010001000000110100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000100011100011110100001011011;
		b = 32'b01100001000110110101111100100011;
		correct = 32'b00000000000100010100100000000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110101100001000010000000000;
		b = 32'b10111101111110001101001000100110;
		correct = 32'b10011100101100001000000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011011000101000001111011101;
		b = 32'b10011110101000101100010101000100;
		correct = 32'b00000010001000101000000101000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000111110000100011011010011;
		b = 32'b00001010111100000110011110101001;
		correct = 32'b00001000111100000100011010000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110111011110100010010001001;
		b = 32'b01011011010011000110101101110100;
		correct = 32'b01001010010011000100000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110101000100011101101001111;
		b = 32'b10010000111000011100101000010000;
		correct = 32'b00010000101000000000101000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111101111001111011010111110;
		b = 32'b01111101010110011001111111100001;
		correct = 32'b01001101000110001001011010100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001001100101100101001010011;
		b = 32'b01110100101100111101001000011100;
		correct = 32'b01110000001100101100001000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010100010001100101000000001;
		b = 32'b10000001111101000010001100100010;
		correct = 32'b00000000100000000000001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100001110001010111101110011;
		b = 32'b00001111000100110010100011110111;
		correct = 32'b00001100000100000010100001110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011000101101100001100101000;
		b = 32'b01011100101010010000100101000100;
		correct = 32'b00011000000000000000000100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011100011110101100000110010;
		b = 32'b00101001011110011110001001000010;
		correct = 32'b00000001000010010100000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111010110100110011101110111;
		b = 32'b11000111101000110101001011111011;
		correct = 32'b00000111000000100100001001110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000000110110011000111000000;
		b = 32'b11111000010000110001010001001101;
		correct = 32'b00011000000000110001000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101001100100011000010001101;
		b = 32'b00110100011000101111111011100001;
		correct = 32'b00100100001000100011000010000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011000001111001110100010011;
		b = 32'b11010001001011110000111111001101;
		correct = 32'b01010001000001110000110100000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110011011101011011001110001;
		b = 32'b10111011101010111110100011001111;
		correct = 32'b10111010001010101010000001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110101010100001010001111010;
		b = 32'b10010001000101010001101001101101;
		correct = 32'b00000000000000000001000001101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110110110111101101110010010;
		b = 32'b10011110011000100111000000101000;
		correct = 32'b10011110010000100101000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111100100000000001111111000;
		b = 32'b00011111000000000011110011000010;
		correct = 32'b00000111000000000000000011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001010011110110011100010110;
		b = 32'b11000000101011001011000011010111;
		correct = 32'b00000000000011000010000000010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110011000100101001101010101;
		b = 32'b10101111101100100111110000010110;
		correct = 32'b00000110001000100101000000010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101011111011010111011000110;
		b = 32'b01100101010001110101111100110111;
		correct = 32'b00000101010001010000111000000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101100111011111011100010101;
		b = 32'b10001010001011101100000100000111;
		correct = 32'b10001000000011001100000100000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100100101010100011010110111;
		b = 32'b00001010111001101100111101111010;
		correct = 32'b00001000100001000100011000110010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000011011110110011110101111;
		b = 32'b00011101111110110001111011110110;
		correct = 32'b00000000011010110000011010100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001110000011101100011110011;
		b = 32'b00001111000001011100011000011010;
		correct = 32'b00000001000000011100000000010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011000010110101001101001000;
		b = 32'b10001111000011110110011110100110;
		correct = 32'b10000011000010110100001100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110001000000000011010101010;
		b = 32'b00110111000110000100010100000100;
		correct = 32'b00010110000000000000010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110111010101101100110110000;
		b = 32'b00000011111011011111000011110101;
		correct = 32'b00000010111010001101000010110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010111001101000101000011111;
		b = 32'b00101010001011101000111101101001;
		correct = 32'b00000010001001101000101000001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001101101001001010111010011;
		b = 32'b10101010111100010100101010111001;
		correct = 32'b00101000101100000000000010010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010010111000000000111000110;
		b = 32'b11001100011001101110001001101100;
		correct = 32'b00001000010001000000000001000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011100000101010100110011100;
		b = 32'b10000010100011010110100011100011;
		correct = 32'b00000010100000000010100010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101101011010001010110011101;
		b = 32'b00001011010100001000100110111000;
		correct = 32'b00000001000000000000000110011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010010010100010011011111101;
		b = 32'b00010010011111000111100001011010;
		correct = 32'b00010010010010000010000001011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101111111100101011010111110;
		b = 32'b00111110001110000111010100111011;
		correct = 32'b00011100001110000101010000111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011110000111111100100010010;
		b = 32'b01100001011010001010001000110100;
		correct = 32'b01100001010000001010000000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001000001010110010010001010;
		b = 32'b01001001010010101110111110010111;
		correct = 32'b00001001000000000110010010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000100111101010001001111101;
		b = 32'b01101101111111010101101010110011;
		correct = 32'b00100000100111000000001000110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010100010011110110011001110;
		b = 32'b10011100000101000001001101100001;
		correct = 32'b10010000000000000000000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010111101110101010000010001;
		b = 32'b00011001010100011010011010101010;
		correct = 32'b00010000010100010000010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000010110011001111011011000;
		b = 32'b10100000101011110001000101110001;
		correct = 32'b00000000000010010001000001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110100110110101100011111100;
		b = 32'b00001000000110000010111110011110;
		correct = 32'b00001000000110000000100010011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101001110001000001011100111;
		b = 32'b00011101100011100010110010001000;
		correct = 32'b00011101000010000000000010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011001010111110011101101010;
		b = 32'b00100111010011001000101101001001;
		correct = 32'b00100011000010001000001101001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010001010100111000101010010;
		b = 32'b11011100010111101011111111111000;
		correct = 32'b01011000000010100011000101010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111111100011111000101111011;
		b = 32'b10000000011001010010110011011100;
		correct = 32'b10000000011000010010000001011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111001101001000101010011001;
		b = 32'b10100100010110010000000111101011;
		correct = 32'b10000100000100000000000010001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010000011101111100100010001;
		b = 32'b11001111110111011111110000110011;
		correct = 32'b11000010000011001111100000010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001000100000011010001111100;
		b = 32'b11001110010111110101100101100011;
		correct = 32'b11000000000100000001000001100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010011100011110111111110011;
		b = 32'b10001001011010000110000111000111;
		correct = 32'b10001000011000000110000111000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011101110100000001101111111;
		b = 32'b11100010011111011100010001000010;
		correct = 32'b00100010001110000000000001000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001111100110110010010001000;
		b = 32'b10011011000101000111011000100100;
		correct = 32'b10011001000100000110010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000010110110111011001011010;
		b = 32'b00011011000011011000011011001100;
		correct = 32'b00010000000010010000011001001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010100110100001000110011111;
		b = 32'b11010001010011000100001010001000;
		correct = 32'b00000000000010000000000010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001100100111101110100110000;
		b = 32'b11101101001010101100100100011000;
		correct = 32'b00000001000000101100100100010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011011100110111100000110101;
		b = 32'b11000000011001000011101110100110;
		correct = 32'b01000000011000000011100000100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100001111011000111011000000;
		b = 32'b01010001111001000110011011011101;
		correct = 32'b00010000001001000000011011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111100101111000100000101101;
		b = 32'b01011010101101010101000110011100;
		correct = 32'b00000010100101010000000000001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000111101101010100000010000;
		b = 32'b00111110000010001010010101001011;
		correct = 32'b00100000000000001010000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011111101110110010111101100;
		b = 32'b01100011110101001001010010111011;
		correct = 32'b01100011110101000000010010101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101111110101011100010111111;
		b = 32'b10101000100100000100101101100100;
		correct = 32'b10001000100100000000100000100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111001100000000111110011100;
		b = 32'b00111111010001000011010100001011;
		correct = 32'b00000111000000000000010100001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111111001110010010000110010;
		b = 32'b10110111010111010111101100100110;
		correct = 32'b00110111010001010010000000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110100111010101100101110101;
		b = 32'b10010011011001011010001100001110;
		correct = 32'b10000010000001010000000100000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001000011001000011101001010;
		b = 32'b10100000010100111101010001111011;
		correct = 32'b10000000000000001000010001001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110000011110100101011010101;
		b = 32'b00101100010100111111001001101001;
		correct = 32'b00101100000000110100001001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110100100011111101101110100;
		b = 32'b01111110100010001110010110110000;
		correct = 32'b01010110100000001110000100110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010010000101101011100100011;
		b = 32'b01101000000111110101000101000011;
		correct = 32'b01000000000000100101000100000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101100101111101001101110111;
		b = 32'b10101000101011010000100000110111;
		correct = 32'b10001000100001010000000000110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111100111010010011001010101;
		b = 32'b10100111101110011110100101010110;
		correct = 32'b10100111100110010010000001010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111100011111011111000110010;
		b = 32'b11011100011011011010011011001001;
		correct = 32'b00011100000011011010011000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111000000011011010010010110;
		b = 32'b11111011111110001010100010111111;
		correct = 32'b10011011000000001010000010010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110000110000010000010001010;
		b = 32'b10100010111110111011011110001100;
		correct = 32'b10000010000110000010000010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011110101101010001011011100;
		b = 32'b00111001001000001101011101010010;
		correct = 32'b00111001000000001000001001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111011011110110101100101010;
		b = 32'b00111110100110011000010000111000;
		correct = 32'b00110110000010010000000000101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101010001110110101111010011;
		b = 32'b00111010101101011101111101001010;
		correct = 32'b00100000000001010100101101000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011001111110000010010001010;
		b = 32'b10000101111001010101000111110011;
		correct = 32'b10000001001001010000000010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000100011011101000011000000;
		b = 32'b00111000100111110111010101111100;
		correct = 32'b00010000100011010101000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110110000010101110101001111;
		b = 32'b11011010101111101101100010001000;
		correct = 32'b00000010100000000101100000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110111010001100010000011001;
		b = 32'b11001111111100010010101001000000;
		correct = 32'b00000110111000000000000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010000000001011000100000100;
		b = 32'b11111011001010110011100010111001;
		correct = 32'b11011010000000000011000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010101010101011011110111101;
		b = 32'b01010111111011110000111101101010;
		correct = 32'b01010010101010100000011100101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010000100110100111110000111;
		b = 32'b10100000000111010001000001010100;
		correct = 32'b10100000000100010000000000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001111110010011101100010111;
		b = 32'b11110000011100110111101010010010;
		correct = 32'b01100000011100010011101000010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001011001110101110100111011;
		b = 32'b00110111000110010110000110001111;
		correct = 32'b00110001000000010100000100001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110001010111101011000011011;
		b = 32'b10010000111101111000001100010111;
		correct = 32'b00000000001000111000001000010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000011010000000001111100100;
		b = 32'b11100111010100101101100100101010;
		correct = 32'b10000000010000000000000100100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110110011001110100001001001;
		b = 32'b01000001110001010010000110011100;
		correct = 32'b00000000110001000010000000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100011100101001100111110101;
		b = 32'b10110010001010100111001100011111;
		correct = 32'b00010000001000100001000100010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011110110101110110101000111;
		b = 32'b10100101011011010010000110000100;
		correct = 32'b10100001010010000010000100000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010101111011001110001101101;
		b = 32'b00000011000101101011011101000100;
		correct = 32'b00000010000101001001010001000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110001011101010101110001001;
		b = 32'b10110011000101100010110011100100;
		correct = 32'b00000010000001100010100010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101010001000011000111100111;
		b = 32'b00100110100101110110010111101000;
		correct = 32'b00100100000001000010000111100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000111100000001000110101100;
		b = 32'b00011010010000001001100010101011;
		correct = 32'b00010000010000000001000010101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000000001001000101110101010;
		b = 32'b11001010000110000010001111010100;
		correct = 32'b11001000000000000000001110000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110011110010111000111111001;
		b = 32'b10011101100101100101000111100110;
		correct = 32'b10011100000100000101000111100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100000100100011100100101011;
		b = 32'b01111011100001111011110010010000;
		correct = 32'b01110000000000100011100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100010100110001110100100110;
		b = 32'b10000100000011001110001111001110;
		correct = 32'b00000100000000000000000100000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001101110000010001001011010;
		b = 32'b11010011000111100011011111010101;
		correct = 32'b00000001000110000010001001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010111111101010010110000010;
		b = 32'b01101011011110100110111101001000;
		correct = 32'b01001010011110100010010100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000111110111101100000001010;
		b = 32'b01011100101110110000011000000001;
		correct = 32'b01001000101110110000000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010100100011100000001000000;
		b = 32'b01001010000010101111010001100011;
		correct = 32'b01001010000000001100000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011101101100010111000100111;
		b = 32'b10000010111011110010010010101010;
		correct = 32'b00000010101001100010010000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011101101101110011000110011;
		b = 32'b11110100011101110010010101001001;
		correct = 32'b00100000001101100010010000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100110000010001100100110110;
		b = 32'b01000000110100001111101111001000;
		correct = 32'b01000000110000000001100100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101011001110111110000100110;
		b = 32'b00010011010100000110001001100000;
		correct = 32'b00000001010000000110000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111000001100111100110011101;
		b = 32'b11001101101111110011011101011001;
		correct = 32'b11000101000001100011000100011001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011011100101011000101110010;
		b = 32'b10111010011100101100111010101011;
		correct = 32'b00011010011100101000000000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101100010001010101101000011;
		b = 32'b00010011000110111110110101001100;
		correct = 32'b00000001000010001010100101000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111010101010110000110011010;
		b = 32'b01011011010000110011110110001000;
		correct = 32'b00010011010000010010000110001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111101100111011100101011111;
		b = 32'b10111111100011010111111100110001;
		correct = 32'b10100111100000010011100100010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100110101101001000011110111;
		b = 32'b01111000110011010011101011011000;
		correct = 32'b00011000110001000001000011010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100111010100001111100101111;
		b = 32'b00011101011001100011011010100110;
		correct = 32'b00010100011000100001011000100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000111000101100011011101100;
		b = 32'b00100000011111000011110010101111;
		correct = 32'b00100000011000000000010010101100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101011011101111100011011011;
		b = 32'b10101000011001001101000100110111;
		correct = 32'b00100000011001001101000000010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011001110111110110001110101;
		b = 32'b10110001000001001000011111000011;
		correct = 32'b00000001000000001000010001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110000101010110000110110001;
		b = 32'b01010000111100010111111111011100;
		correct = 32'b00000000000100010110000110010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001101011000110111100110101000;
		b = 32'b01101101010100101010000000000010;
		correct = 32'b00001101010000100010000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111011010001111101010101000;
		b = 32'b00101100011000110000101100101000;
		correct = 32'b00100100011000000000101000101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100110001111101001000111011;
		b = 32'b00001111100100010100011100001001;
		correct = 32'b00001100100000010100001000001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000101011110000001011001111;
		b = 32'b00110011010001000001100011101011;
		correct = 32'b00100000000001000000000011001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000000011010010000010101101;
		b = 32'b10111101100110000110011011110011;
		correct = 32'b00110000000010000010000010100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000001001110000101110101000;
		b = 32'b11011001000110010000011010100001;
		correct = 32'b10011000000000010000001010100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100011001000001001011001110;
		b = 32'b10100001001101110111001111010000;
		correct = 32'b10000000001001000001001011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110111011100101000010101010;
		b = 32'b00001111110001110011101001011110;
		correct = 32'b00001110110001100001000000001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100001011111001111111010100;
		b = 32'b00100001110011010110001011000101;
		correct = 32'b00100000000011010000001011000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001010101100111000111110111;
		b = 32'b00000000010011000101101101010001;
		correct = 32'b00000000010001000101000101010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010100000100010101001010001;
		b = 32'b11110100110000101111011000111000;
		correct = 32'b00000000100000100010001000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110010000001000011110010101;
		b = 32'b10111101011100011110010100111111;
		correct = 32'b10001100010000001000010100010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110000111000100111110010000;
		b = 32'b11001100001110000010000010110001;
		correct = 32'b00000100000110000000000010010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011000001110111110111110000;
		b = 32'b00100011011011100000100010111100;
		correct = 32'b00000011000001100000100010110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010011111101111000111110010;
		b = 32'b10100100011111101011110001110000;
		correct = 32'b10000000011111101011000001110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001101011001111110101011001;
		b = 32'b00110111111001111100001011111010;
		correct = 32'b00000001101001001100000001011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001001001000010100001011100;
		b = 32'b11000001001011111111010101111001;
		correct = 32'b01000001001001000010000001011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110001010101110001011000001;
		b = 32'b00110001001101000100110111000110;
		correct = 32'b00100000001000000100000011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101111010111011011110011010;
		b = 32'b00111101110111100011011010001001;
		correct = 32'b00111101110010100011011010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011100000000111100110000000;
		b = 32'b00111110011001101001101010110001;
		correct = 32'b00101010000000000001100010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000011010010011101111010001;
		b = 32'b01101101010000110011110000010001;
		correct = 32'b00100000010000010011100000010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100000010101100011110110100;
		b = 32'b01000001110001000000111101000001;
		correct = 32'b01000000000000000000011100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010010011011000100111001111;
		b = 32'b00011100000000011110011001010110;
		correct = 32'b00000000000000011000000001000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100000100111111111111111001;
		b = 32'b00110000111001000010110100000000;
		correct = 32'b00100000000000000010110100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111100011001010011111010100;
		b = 32'b00110011001010100100011001000001;
		correct = 32'b00000011000010000000011001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111101010010001010100100111;
		b = 32'b01101011001110011001001001000101;
		correct = 32'b01000011001010010001000000000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010100110111111010111100000;
		b = 32'b01100110011111111100100111101110;
		correct = 32'b01000010000110111100000111100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001110010111010110111100000;
		b = 32'b00010100111111100100101001011000;
		correct = 32'b00000000110010100000100001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110000011110110101000001101;
		b = 32'b01011100110100101101101011111000;
		correct = 32'b01011100000000100100101000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000101010100010001101010011;
		b = 32'b10111001111011110110001111100001;
		correct = 32'b10110000101010100010001101000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000001011001010001011111011;
		b = 32'b11000110111000101110011101110111;
		correct = 32'b11000000001000001010001001110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101001101000010000110011010;
		b = 32'b01110001100010011111101000110010;
		correct = 32'b01110001000000000010000000010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010100101110101110000001010;
		b = 32'b10011100010001011010110000110001;
		correct = 32'b00010000000001010000110000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010111001001101111001011010;
		b = 32'b11000110100000010011010011110000;
		correct = 32'b01000010100000000001010001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110101110000011101011011001;
		b = 32'b11110000011010100111001110111110;
		correct = 32'b01010000001010000011001010011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001000000011110001010000110;
		b = 32'b10001100100100000110101110010100;
		correct = 32'b10001000000000000110001010000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011101011101111000011101000;
		b = 32'b00010101011001111101100011010100;
		correct = 32'b00000001001001101101000011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100100111001000111110100010;
		b = 32'b10111001001101011111101110111000;
		correct = 32'b00100000000101001000101110100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011001000010101001011001010;
		b = 32'b01000101110101011000001110100010;
		correct = 32'b00000001000000010000001010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100111001001110100111101111;
		b = 32'b00000011101001011001101101110010;
		correct = 32'b00000000101001001000100101100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011000010011110011010010001;
		b = 32'b10010101010010101110111011100010;
		correct = 32'b10000001000010001110011010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001010111011101101101000111;
		b = 32'b00001100000000100000011010111100;
		correct = 32'b00001000000000000000001000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111000000111110111101010111011;
		b = 32'b10000111010110111010111001011100;
		correct = 32'b00000000000110110010101000011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010001010111111111100010010;
		b = 32'b01011100110100001110111010010000;
		correct = 32'b01000000000000001110111000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001010100100010001101110101;
		b = 32'b00000010011110000001011110011100;
		correct = 32'b00000000010100000000001100010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000011010001000111000011000;
		b = 32'b00101011000101101011010001111111;
		correct = 32'b00001000000000001000010000011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111010110100001000011001100;
		b = 32'b01011101010010101101001110101110;
		correct = 32'b01001101010010100001000010001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000000001001011011000100101;
		b = 32'b10000011110111011000010000001010;
		correct = 32'b00000000000001001000010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000000111111011100001100001;
		b = 32'b00001000111001000101110101110110;
		correct = 32'b00000000000001000001100001100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100011111001011000011010001;
		b = 32'b10010001111100101101011011110101;
		correct = 32'b00010000011100001001000011010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111111000001110001010101101;
		b = 32'b01100001110111110011010010011010;
		correct = 32'b00000001110000000010000010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001010100101111110011101111;
		b = 32'b01010000110000110011111000000110;
		correct = 32'b01000000010000100011110000000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111100101101010010011101100;
		b = 32'b01100010011100110111010001110111;
		correct = 32'b00100010000100100010010001100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000111010110011101001100110;
		b = 32'b11100101011001010000111100101011;
		correct = 32'b10100000011000010000101000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000100100111000001011100110;
		b = 32'b00101001101011010001111010010011;
		correct = 32'b00001000100000010000001010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011110010101111100111001101;
		b = 32'b11101100011110111011111110100000;
		correct = 32'b11000000010010101011100110000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010010011001001000100101000;
		b = 32'b11000101010000101110110101011110;
		correct = 32'b11000000010000001000000100001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101111111111010000101001110;
		b = 32'b11101010110111010010001001111000;
		correct = 32'b11100000110111010010000001001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011100100000011111111001011;
		b = 32'b11100000001111100100110101010101;
		correct = 32'b01000000000100000000110101000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100101001011111001011100000;
		b = 32'b10011010010110000100001010100100;
		correct = 32'b00010000000000000100001010100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001010010010100100000110101;
		b = 32'b01100100111001001010011110000001;
		correct = 32'b01100000010000000000000000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000001110000110111100010011;
		b = 32'b11110010111110011110110011001000;
		correct = 32'b01110000001110000110110000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111000101101000100111011100;
		b = 32'b01000000011001011010010001001011;
		correct = 32'b01000000000001001000000001001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001110100000000000011000000;
		b = 32'b01100010101111010110001001001101;
		correct = 32'b01000000100100000000000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000101011100001010111101011;
		b = 32'b00101001010100110001001111111110;
		correct = 32'b00101000000000100001000111101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100101111110101100010000010;
		b = 32'b01010110011111001101001010110001;
		correct = 32'b01010100001111000101000010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011010001011000110010111111;
		b = 32'b01111000010100010010011000010101;
		correct = 32'b01001000010000010000010000010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100110010100000111101111010;
		b = 32'b11001010000110110111001101101011;
		correct = 32'b01000000000010100000001101101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101100110001101011100011010;
		b = 32'b11101111000100100110001111001000;
		correct = 32'b01101101000100000100001100001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110111110000110011110101100;
		b = 32'b01010110000101100101011000110111;
		correct = 32'b00000110000100000100011000100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110110101011100010011110000;
		b = 32'b10011011010101110000010000000111;
		correct = 32'b10011010010101010000010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111000000001011100111110011;
		b = 32'b00111011000010001000011000111101;
		correct = 32'b00011011000000001000000000110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111010010010101110010011101;
		b = 32'b01101000010011111110011011100010;
		correct = 32'b01001000010010010100010010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001100011101110100101000000;
		b = 32'b11010010010001010110100001111101;
		correct = 32'b00000000000001000110100001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000011101100001010101101111;
		b = 32'b10110001011111100100000000100110;
		correct = 32'b00000000011101100000000000100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100000001010000110001111011;
		b = 32'b11001011001110000001001110101010;
		correct = 32'b00001000000000000000000000101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110001001011100010111110001;
		b = 32'b01101110001011100011101001111111;
		correct = 32'b00101110001001000000000001110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001101001100101010010011111;
		b = 32'b11011101100100110001101010111110;
		correct = 32'b11000001100000100001000010011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100010101111000110000010000;
		b = 32'b01100101101011111100010000110111;
		correct = 32'b00000100000001111000010000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010011100001100010101110101;
		b = 32'b01011100110001101010011000001100;
		correct = 32'b00001000010000001000010000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110110001110111010011010110;
		b = 32'b01010001001000001001110000000111;
		correct = 32'b01000000000000000001010000000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011001000111110101011011011;
		b = 32'b11101100101101101000010101000101;
		correct = 32'b00000000001000101000000001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011100000100010110001110011;
		b = 32'b01110001000010010010111010111101;
		correct = 32'b01110001000000000010110000110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101100011110000101111001110;
		b = 32'b11001110000101111100101010011010;
		correct = 32'b01000100000001110000101010001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000101111010011100101011011;
		b = 32'b00100100110111011111110111101100;
		correct = 32'b00100000100111010011100101001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010110001000100110011100000;
		b = 32'b00001101100000001100110000011101;
		correct = 32'b00000000100000000100110000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010111000011001100010011110;
		b = 32'b10011000100110111111001100110001;
		correct = 32'b00011000100000011001000000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011101111001000100001100101;
		b = 32'b10010101000001011000101010001010;
		correct = 32'b10000001000001001000100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111110100110011111010000010;
		b = 32'b11001000100000011101001110111111;
		correct = 32'b01000000100000010001001010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001101001101100101111111011;
		b = 32'b10110100110101101010011100010111;
		correct = 32'b00110000100001101000001100010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100100111100111010111110011;
		b = 32'b00000010100011011001001010111100;
		correct = 32'b00000000100011000001000010110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111011111011111010000100110;
		b = 32'b11000101011000111100100100101111;
		correct = 32'b10000101011000011100000000100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111111100100111001010000111;
		b = 32'b01101010001000101100011011010101;
		correct = 32'b00100010001000100100001010000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000101000101011010101110111;
		b = 32'b10010111100001001110000101100110;
		correct = 32'b10000000100000001010000101100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000101010010101001011100101;
		b = 32'b11101110101101100110101110110001;
		correct = 32'b11001000101000000100001010100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011001111000001011100110011;
		b = 32'b11101010101000110111001111100001;
		correct = 32'b11100010001000000001001100100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011101000010100111010000000;
		b = 32'b00010001010101001010011100001011;
		correct = 32'b00000001000000000000011000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101100100110010010000000101;
		b = 32'b10011001101110110111001011101010;
		correct = 32'b10011001100100110010000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100000010001100100010001101;
		b = 32'b00101000110100110011101110010011;
		correct = 32'b00101000000000000000100010000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001001110000000110001010111;
		b = 32'b01000001001100011110111111000011;
		correct = 32'b01000001001100000000110001000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100000100000110101010000010;
		b = 32'b10111100010001001000100001010101;
		correct = 32'b00111100000000000000100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100111101110101111010110111;
		b = 32'b00100110111100111110011101010111;
		correct = 32'b00000100111100110100011000010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000001100011001011001100000;
		b = 32'b01011110100111000101111110000111;
		correct = 32'b01000000000100000001011000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011101000000110010101100100;
		b = 32'b00010000100010010100000110100110;
		correct = 32'b00000000100000000100000100100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101101111000000001101110100;
		b = 32'b11101010011010111001101010001100;
		correct = 32'b10101000001010000000001000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011110000100011011101101010;
		b = 32'b10110001100101001010001011111101;
		correct = 32'b10110001100000000010001001101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101001011011011110011100101;
		b = 32'b01001011011000011010100011010110;
		correct = 32'b00000001001000011010100011000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100011111010100011110000111;
		b = 32'b10010100000011101100110000011111;
		correct = 32'b00010100000011000100010000000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110111101101101101110100000;
		b = 32'b00010011010000000101001101111100;
		correct = 32'b00000010010000000101001100100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011101001101010001010111111;
		b = 32'b00100100011010001100110110010001;
		correct = 32'b00100000001000001000000010010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111000100100000101111111111;
		b = 32'b10100001001001101111111010001111;
		correct = 32'b00100001000000100000101010001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001110100111100111011111011;
		b = 32'b00010001101010101001010000011111;
		correct = 32'b00000001100000101000010000011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011111010000000010100110011;
		b = 32'b11100011011100111101011111001000;
		correct = 32'b00000011011000000000010100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111110101100000110100101000;
		b = 32'b01100101111001001111100110111111;
		correct = 32'b00000101110001000000100100101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011010110011100001100111000;
		b = 32'b10110011101001011010010111000000;
		correct = 32'b00000011000000011000000100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101111000111001110011111100;
		b = 32'b00110111000110000101101110001000;
		correct = 32'b00000101000000000001100010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011011100100101101100111101;
		b = 32'b10101101001001111110111010001010;
		correct = 32'b00100001001000100100101000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011110000111011110101010011;
		b = 32'b01011001001110111111100011111110;
		correct = 32'b01000001000000111011100001010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011011100100100100001111111;
		b = 32'b10000111100101110100110001101011;
		correct = 32'b10000011000100100100100001101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011000011100001000100110001;
		b = 32'b10100000101001111111001110111101;
		correct = 32'b00100000000001100001000100110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000111001111011111001110111;
		b = 32'b11100101010000000000100010010101;
		correct = 32'b11100000010000000000100000010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000000110111110010100011000;
		b = 32'b01010111110011111100001111100011;
		correct = 32'b00010000000010111100000100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001110110001110111001101000;
		b = 32'b11010101111101101101010010110000;
		correct = 32'b01000001110100001100010000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111010111100111010000101000;
		b = 32'b01011011010100110011011101010110;
		correct = 32'b00001011010100100011010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101000110011010100010010000;
		b = 32'b10110111011101111001110110111101;
		correct = 32'b00110101000100011000100010010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100001101011001101001110000;
		b = 32'b01010101110001010001000011010110;
		correct = 32'b00010100000001010001000001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011001001111001010001001001;
		b = 32'b11111001101010001101000101110000;
		correct = 32'b00100001001000001001000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011100010110010001110001000;
		b = 32'b00010111111100010010110100111100;
		correct = 32'b00000011100000010010000100001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010011011101011100000100011;
		b = 32'b10100111001101011010111101111010;
		correct = 32'b00000010001001001010100000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010100111110000101001011110;
		b = 32'b01100100011101101001010011011111;
		correct = 32'b00000000000101100000000001011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011011101001010100111111011;
		b = 32'b01101110111001001001000100111110;
		correct = 32'b01001010011001001000000100111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100111101100111101001011010;
		b = 32'b00000001010000111100010111100111;
		correct = 32'b00000000010000100100000001000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101100101000000010001010010;
		b = 32'b10011010110000000101111111011101;
		correct = 32'b10011000100000000000010001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001010100010011011111101001;
		b = 32'b01110100101001100000001100110000;
		correct = 32'b00100000000000000000001100100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100101110101101111111111110;
		b = 32'b00110000110000000101111101010000;
		correct = 32'b00100000100000000101111101010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000010111011101011101101011;
		b = 32'b10100000010110111110000111010110;
		correct = 32'b10100000010110011100000101000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101001011010111100011111100;
		b = 32'b11010011000100010111110000010010;
		correct = 32'b11010001000000010111100000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010111111000001100101100001;
		b = 32'b11110010101101001011110011010010;
		correct = 32'b01100010101101000001100001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010001110110011000001000000;
		b = 32'b11101110111011101011000001000111;
		correct = 32'b01000010001010100011000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000100010010000100101011110;
		b = 32'b11001010100111100011100011001011;
		correct = 32'b11001000100010000000100001001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001110000001111100011110000;
		b = 32'b00101010010010000001010000100100;
		correct = 32'b00000000010000000001000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111001110111100111001010001;
		b = 32'b01111011011111111110011011111011;
		correct = 32'b00110011001110111100011001010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011110000000000001001001001;
		b = 32'b10011001001000001010000110110000;
		correct = 32'b10000001000000000000000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101011101011000101100011000;
		b = 32'b01010101011000111100010100101110;
		correct = 32'b01000101011000011000000100001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000100000001010111100001111;
		b = 32'b00110110110001001110011010010000;
		correct = 32'b00010000100000001010011000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011101001110110000000010001;
		b = 32'b00110101001011001000111010000011;
		correct = 32'b00110001001001000000000000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111100010101110010000100101;
		b = 32'b01011001101111111001111000111110;
		correct = 32'b01001001100010101000010000100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000011001001100010111101010;
		b = 32'b00110011010110100111010011000100;
		correct = 32'b00010000010000000100010011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100010011010011000011101100;
		b = 32'b11001100111100100011001111000111;
		correct = 32'b00000100010000000011000011000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100100011001110100011101010;
		b = 32'b00100101000111111101000110010111;
		correct = 32'b00100100000011001100000010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011111111100011001010011101;
		b = 32'b11000011101111110001101101110011;
		correct = 32'b10000011101111100001001000010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110101100000011011010001001;
		b = 32'b00001101101011010110110110100101;
		correct = 32'b00001100101000000010010010000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001100111010001110100101100;
		b = 32'b00011111010000110001010110010010;
		correct = 32'b00000001000000010001010100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001000010011011001101111111;
		b = 32'b11000000111111000000110111010111;
		correct = 32'b11000000000010000000000101010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001011010101100000110011000;
		b = 32'b11100000101010100001100010011110;
		correct = 32'b11000000001010100000000010011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100011100000110100011011001;
		b = 32'b10001011010100110001100001011000;
		correct = 32'b10000000010100000000100001011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110101001001010001001100010;
		b = 32'b10010101100110100010011001111110;
		correct = 32'b10010100100000000010001001100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011110110011110100001000010;
		b = 32'b10011011111110111010101100100100;
		correct = 32'b00000011110110011010100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111001100110010000011010000;
		b = 32'b11010001001011100101100011101100;
		correct = 32'b10010001001000100000000011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110101001100001010111001011;
		b = 32'b00000011101110100101111101000111;
		correct = 32'b00000010101000100001010101000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101011101001010101111011000;
		b = 32'b00110011000110101110011001100010;
		correct = 32'b00100001000100001010001001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010101010100101110101110111;
		b = 32'b10100111101000000111101010111100;
		correct = 32'b00000010101000000101100000110100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100011101011011111101110011;
		b = 32'b11101010000101111010010011000010;
		correct = 32'b00001000000101011010010001000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101111001010101010001000100;
		b = 32'b00010001000001110001010111000011;
		correct = 32'b00010001000001010001010001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111001011000011100000001111;
		b = 32'b11010101101110111010011001100100;
		correct = 32'b01000101001010000010000000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101001011001101001101000100;
		b = 32'b10101110100001101100100110110111;
		correct = 32'b10100100000001001100000100000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011011111010001011000111001;
		b = 32'b10101001000101011011101011000001;
		correct = 32'b10000001000101010001001000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111011100110110011000010101;
		b = 32'b10001110001010010101001010100011;
		correct = 32'b00000110001000010100001000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111101000110000110110111011;
		b = 32'b00100101101010111000001111101011;
		correct = 32'b00000101101000110000000110101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111011110001110001000001100;
		b = 32'b01100110000000011000001000000010;
		correct = 32'b00000110000000001000001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010010010000111110110111000;
		b = 32'b01001000100110110011101101101001;
		correct = 32'b00001000000010000011100100101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101101011101100011111000101;
		b = 32'b00100001011101011011110100000111;
		correct = 32'b00100001001001001000010100000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000110001101010000010011000;
		b = 32'b11011011100111001111100110000111;
		correct = 32'b11010000100001001010000010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111001011100100110010000000;
		b = 32'b11100010000100010110001001000000;
		correct = 32'b00100010000000000100000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011101100010101111001010010;
		b = 32'b11101001001010000000110110000111;
		correct = 32'b01001001001000000000110000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111111101010111001101110101;
		b = 32'b01001011111111000111100011000001;
		correct = 32'b00000011111101000111000001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010111000110011110010101110;
		b = 32'b11110001000011001011111111010000;
		correct = 32'b01000000000000000011110010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100000111000010011011011011;
		b = 32'b01111101010101100010111000100111;
		correct = 32'b01010100000101000010011000000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111100001010010010000111111;
		b = 32'b01110110000101101010000000001010;
		correct = 32'b01010110000001000010000000001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111011000110010001110100110;
		b = 32'b10001001001011011010101111000101;
		correct = 32'b10000001001000010010001110000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110001010101111111011001000;
		b = 32'b01111000111011101001100111101000;
		correct = 32'b01000000001010101001100011001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100110101001101100100111010;
		b = 32'b01011000000010010111101000110110;
		correct = 32'b01011000000000000101100000110010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111101111000011110100010001;
		b = 32'b00010010000111000000000101000110;
		correct = 32'b00000010000111000000000100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110110001101110111010100100;
		b = 32'b11011001000000011100101000111101;
		correct = 32'b10010000000000001100101000100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101011010101010001110100011;
		b = 32'b11001111100001011110111000100001;
		correct = 32'b10001101000000001010001000100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000001100011110010010100011;
		b = 32'b10000101100010000110101001101100;
		correct = 32'b10000000000000000110000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011001111111011010110011110;
		b = 32'b00101110111101010011110001100110;
		correct = 32'b00000010001101010011010000000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110111100110100100101111010;
		b = 32'b00111001001111001110010010011010;
		correct = 32'b00000000001100000100000000011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101000010001101010000010110;
		b = 32'b10010011010000010100101110100000;
		correct = 32'b00010001000000000100000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101101111001100010111101100;
		b = 32'b00000111001010001001000010011001;
		correct = 32'b00000101001010001000000010001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010101100100000011000110110;
		b = 32'b00000011001100011011110100101001;
		correct = 32'b00000010001100000000010000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000100110101110011011001110;
		b = 32'b00100110111001101010010001110100;
		correct = 32'b00000000100000101010010001000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010100011010011110101000010;
		b = 32'b11011111101111001001000000101100;
		correct = 32'b11001010100011000001000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110010111011011010100010001;
		b = 32'b11000010000100011011101001111100;
		correct = 32'b00000010000100011011000000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001111010101000100010011001;
		b = 32'b10000000001000111110011011011001;
		correct = 32'b10000000001000101000000010011001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010111110010000010111101001;
		b = 32'b01110011110001010010001101010100;
		correct = 32'b00010010110000010000000101000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010011101000101001110101000;
		b = 32'b00100101101110110011010110010011;
		correct = 32'b00000000001100000001000110000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101110010101001100101111110;
		b = 32'b11110110100110001101001100101000;
		correct = 32'b01010100100010001001000100101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010100101110010001101101010;
		b = 32'b01001010101000011011010101011000;
		correct = 32'b00000010100000010010000101001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011111111101100010101010000;
		b = 32'b01000101000000100001010011100000;
		correct = 32'b01000001000000100000010001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001111000111011000110111110;
		b = 32'b11010001001111010011111000011101;
		correct = 32'b01000001001000010011000000011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011101000101100000101001100;
		b = 32'b01101101111110000100011101110110;
		correct = 32'b01101001101000000100000101000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010110101100011000001110011;
		b = 32'b01010010101101001110101010001001;
		correct = 32'b00000010100101000010000000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110010111101100001001001011;
		b = 32'b01011001011110000000010111101011;
		correct = 32'b00001000010110000000000001001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110000011100100010010010010;
		b = 32'b11110001011000101101100110110001;
		correct = 32'b10010000000000100100000010010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110111000011110000111001111;
		b = 32'b01100001100110010101110000110111;
		correct = 32'b01100000100000010100000000000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110000000111001011011111010;
		b = 32'b10110111000011100011100101110101;
		correct = 32'b10110110000000100001000001110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000101101100001010001011111;
		b = 32'b01100000011000010001110111110111;
		correct = 32'b00000000001000000001010001010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111010110100101001001011101011;
		b = 32'b00111101010011101100010110010011;
		correct = 32'b00111000010000101000000010000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101010000000100000100000010;
		b = 32'b00000000110111111111010111111110;
		correct = 32'b00000000010000000100000100000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110010010111111101010010001;
		b = 32'b10011111010001011100001110100010;
		correct = 32'b00001110010000011100001010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100001001100001101001010101;
		b = 32'b10111101010100000010010110011100;
		correct = 32'b00100100000000000000000000010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010100011101010010101001100;
		b = 32'b10100110000101101101011001111110;
		correct = 32'b00100010000001101000010001001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001111001010101011111000001;
		b = 32'b01011110000011111001111101101010;
		correct = 32'b00000000000001010001011101000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110111001100000101011001001;
		b = 32'b00110011010011111101011011010101;
		correct = 32'b00110010010001100000001011000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101000101101001100001010100;
		b = 32'b11110001100010110110011010110111;
		correct = 32'b01100001000000100000000000010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011100111011001111101001000;
		b = 32'b00111001100001001001101110100100;
		correct = 32'b00001001100001001001101100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101001010000100100011101111;
		b = 32'b11010111101110110000101001100110;
		correct = 32'b11000101001010000000100001100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010101100111011011100110111;
		b = 32'b01100000011110001110110100000101;
		correct = 32'b00100000001100001010010100000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000010010100001111010100111;
		b = 32'b00111101110111111011010011010101;
		correct = 32'b00011000010010100001010010000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111111100001101111111001001;
		b = 32'b11011111001001010010011101000000;
		correct = 32'b10001111001000000000011101000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100111000001110110011000101;
		b = 32'b01100000111001000100110111101000;
		correct = 32'b01000000111000000100110011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100010110000100001001110100;
		b = 32'b01101000100100010001010111101000;
		correct = 32'b01100000000100000000000001100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010001110000010011100111101;
		b = 32'b00100110100111110011000111000011;
		correct = 32'b00100010000110000010000100000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100010101110110100010010001;
		b = 32'b01010101111010011010010000011101;
		correct = 32'b00010100010000010010000000010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000001111001001001110000000;
		b = 32'b00001000000110011101111000111000;
		correct = 32'b00001000000110001001001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110101100001011111111010001;
		b = 32'b01010001011111111001111101111001;
		correct = 32'b01000000001100001001111101010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010011001111110101011101001;
		b = 32'b01010010001110000011011111011110;
		correct = 32'b01010010001000000010001011001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110101010001010110110100001;
		b = 32'b00101010001100110011001011100001;
		correct = 32'b00101010001000000010000010100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011101011001000010111110110;
		b = 32'b10101000010100111110001110000100;
		correct = 32'b10001000000000001000000110000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011111110001001001110001010;
		b = 32'b10001100101011001110011001100100;
		correct = 32'b00001000101010001000001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000000011011111001100010001;
		b = 32'b00011000010011001111011001010100;
		correct = 32'b00001000000011001111001000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111010000001010111110111000;
		b = 32'b00111111011110111110100100011010;
		correct = 32'b00001111010000001010100100011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111101011001110001101001101;
		b = 32'b00010011001101010000100111010101;
		correct = 32'b00000011001001000000000101000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100101101011100011100010111;
		b = 32'b11001110111110111101001000001110;
		correct = 32'b01001100101100011100001000000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110110010011101110011000110;
		b = 32'b11001101010000010011100001100011;
		correct = 32'b01001100010000010001100001000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101101110011001001100001110010;
		b = 32'b10110010110010100101000111011001;
		correct = 32'b00100000110010000001000001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110111010011010111001000100;
		b = 32'b00001001000001100010101101000111;
		correct = 32'b00001000000000000010101001000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100100001011101110010001100;
		b = 32'b00101001100011101111111011110010;
		correct = 32'b00100000100001001101110010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010001000010100010010011000;
		b = 32'b01100001001111111011001100001101;
		correct = 32'b01100000001000010000000000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001101110010100010001010110;
		b = 32'b00111000101000011111000010100001;
		correct = 32'b00110000101000010100000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111111110101001000000000000;
		b = 32'b00100000001100100110001110110100;
		correct = 32'b00000000001100100000000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000010001111110010100001101;
		b = 32'b10011100100011101111011010001111;
		correct = 32'b10000000000001101110010000001101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111011010011100101100101011;
		b = 32'b01110001001011010001110000011010;
		correct = 32'b01100001001010010000100000001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001111110100010001100111110;
		b = 32'b00101110000100101101100000100010;
		correct = 32'b00100000000100100000000000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011011000100000011001000001;
		b = 32'b10001001110000001001110100111101;
		correct = 32'b10000001010000000000010000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010011110100100111111000011;
		b = 32'b01011011111001111000110101100010;
		correct = 32'b00011010011000100000110101000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001110011100001101011100100;
		b = 32'b00010001011010011010001101010110;
		correct = 32'b00000001010010000000001001000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000100001011011010110100101;
		b = 32'b10101011101111001010100101110000;
		correct = 32'b00100000100001001010000100100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100001100101010010101100101;
		b = 32'b01001001101110110010001110100100;
		correct = 32'b00000000001100100010000100100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010010011000001010001011010;
		b = 32'b00101101001101100100101111111101;
		correct = 32'b00000000000001000000000001011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111011011111001000111110110;
		b = 32'b10000111111101110110000010011110;
		correct = 32'b00000111011001110000000010010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100001011111001001001100110;
		b = 32'b11001010010010110110000010111000;
		correct = 32'b00001000000010110000000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001000001111010010001000000;
		b = 32'b11100010001000101101110110001001;
		correct = 32'b11100000000000101000010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000010110000010110100110100001;
		b = 32'b00110010010001001101100010101110;
		correct = 32'b00000010010000000100100010100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011001001111000111001001101;
		b = 32'b00011111110000011111101100101000;
		correct = 32'b00011011000000011000101000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101011000110101010000000100;
		b = 32'b11010101110111111011101101010110;
		correct = 32'b10010101010000110001000000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101011011101000100101011100;
		b = 32'b10110011101000000001011100101110;
		correct = 32'b10100001001000000000000100001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110101011001010001111101000;
		b = 32'b01101111100011101010001110010110;
		correct = 32'b00101110100011001010001110000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011011100011000011110101010;
		b = 32'b00001101010100000000101110111000;
		correct = 32'b00001001010100000000001110101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111101011101111100100001101;
		b = 32'b00110100001010100000110110010001;
		correct = 32'b00010100001010100000100100000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101111111111100111110101101;
		b = 32'b10000011001001111110000101100110;
		correct = 32'b00000001001001111100000100100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100111110010011111000101110;
		b = 32'b10000001101110110010001100101110;
		correct = 32'b00000000101110010010001000101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001010001000111001010001111;
		b = 32'b11100110010001101100000010101010;
		correct = 32'b11100000010001000100000010001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101111110000000100111110111;
		b = 32'b00111101011011100101101110011111;
		correct = 32'b00101101011010000000100110010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100110001111101000110010110;
		b = 32'b10000010011100001001100111111100;
		correct = 32'b00000000010000001001000110010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010100011110111011110000001;
		b = 32'b10101111000011001110101101111000;
		correct = 32'b00101010000011000110001100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100011001111011011111101000;
		b = 32'b10110101101011000111010110110100;
		correct = 32'b00100100001001000011010110100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110110100111101000001000100;
		b = 32'b10011110111001000001110000001101;
		correct = 32'b00010110110000000001000000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100010010001011001111010001;
		b = 32'b00010101111001110000001101110011;
		correct = 32'b00000100010000000000001101010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001100110011001101001001101;
		b = 32'b01010001010010001001000111001101;
		correct = 32'b00000001000010001001000001001101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111011010010010010011000101;
		b = 32'b00011110001001011110000000100100;
		correct = 32'b00000110001000010010000000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010101001111010101101100011;
		b = 32'b11111111111110011000000000110011;
		correct = 32'b00111010101000011000000000100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010000011100000110111111001;
		b = 32'b01101100110001110110011011101100;
		correct = 32'b00100000000001100000010011101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100010000101111110100100011;
		b = 32'b01100101001001001011001100011111;
		correct = 32'b00000100000000001011000100000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010011101100000001101111001;
		b = 32'b11011100110111111011101100010010;
		correct = 32'b11001000010101100000001100010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111010011100010011010011100;
		b = 32'b01100010101100110111011110011001;
		correct = 32'b01000010000000100010011010011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011010101111010100110111110;
		b = 32'b00100110110000001100000110000000;
		correct = 32'b00000010010000001000000110000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100011000110000111011010101;
		b = 32'b10011100110100001110010101000011;
		correct = 32'b00011100010000000000010001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111000000000101110110110010;
		b = 32'b11011001011010010110101101111101;
		correct = 32'b11000001000000000100100100110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001000100011101011010011100;
		b = 32'b00001100001110100000001110111000;
		correct = 32'b00000000000100000000001010011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000010011010011011011000101;
		b = 32'b00111110100010010001101110001100;
		correct = 32'b00101000000010010001001010000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111111101111000100110000011;
		b = 32'b01111011110000111010010100010110;
		correct = 32'b01011011110000111000000100000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110001111000001110111001110;
		b = 32'b01010101101011101001000110010000;
		correct = 32'b01000100001011000001000110000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111010000101000110100110000;
		b = 32'b11100001001101111101011001001011;
		correct = 32'b11000001000000101000010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011011101101001100000000111;
		b = 32'b01000001101001000000110000001000;
		correct = 32'b01000001001001000000100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111000110000011110110111111;
		b = 32'b10001001011001001000000010000000;
		correct = 32'b00001001000000000000000010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000110100011110010110010110;
		b = 32'b10100111111101010000101110001011;
		correct = 32'b10100000110100010000000110000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000111000011000001101100001;
		b = 32'b01101111101111110111000101110010;
		correct = 32'b00001000101000010000000101100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000100101101000001011100111010;
		b = 32'b00101000000000110110010110101100;
		correct = 32'b00000000000000000000010100101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100001111111000010100011101;
		b = 32'b00010011010110111100100110010100;
		correct = 32'b00010000000110111000000100010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111101101100010011010101110;
		b = 32'b11001111111111110111100111110001;
		correct = 32'b10001111101101100010000010100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111010000010011111001100101011;
		b = 32'b11000110001011111110011110100110;
		correct = 32'b11000010000010011110001100100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001011001101110110011011110;
		b = 32'b01011111111000001111110001100100;
		correct = 32'b00000001011000001110110001000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011101101101100010001110101;
		b = 32'b00011000100000111100000101111100;
		correct = 32'b00010000100000101100000001110100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111000100100111001111101110;
		b = 32'b01111111111101111100011101110001;
		correct = 32'b00101111000100100100001101100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111100010010101001100010011;
		b = 32'b11001111011100100000011101100101;
		correct = 32'b11000111000000000000001100000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001101111010100101100101001111;
		b = 32'b11011011011101101111010011001011;
		correct = 32'b00001001011000100101000001001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101001110010110111110100100;
		b = 32'b11000000100001111010010001000100;
		correct = 32'b10000000000000010010010000000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011011100001011110001100101;
		b = 32'b00000101010000010100111101111110;
		correct = 32'b00000001010000000000110001100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111011110000000011001011111;
		b = 32'b10001100011110001000110110111111;
		correct = 32'b10001100011110000000010000011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100001011100101001001000101;
		b = 32'b01010001011000001111111101011011;
		correct = 32'b01010000001000000101001001000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110100111010011001100001100;
		b = 32'b01111101110111110101001111101101;
		correct = 32'b00000100100111010001001100001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100011011110000110000001101;
		b = 32'b00011101010100011011010000101001;
		correct = 32'b00000100010000010000010000001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100000111100110101101001110;
		b = 32'b10111111100001110011001110010000;
		correct = 32'b00011100000001100010001100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000110110111110011001011011;
		b = 32'b10000111001111100000110101001111;
		correct = 32'b00000000000110100000010001001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001001001011101111001110110;
		b = 32'b01101010101111011001100001100011;
		correct = 32'b00001000001001011001100001100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000110100000001111010111010;
		b = 32'b00011000100010110011000111100010;
		correct = 32'b00010000100000000001000010100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101001000011111011111000001;
		b = 32'b10111001110001100001011111100110;
		correct = 32'b00011001000000000001011111000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110100001000011100000010011;
		b = 32'b10001001101000000110000010001001;
		correct = 32'b10001000100000000010000000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101011000110001100011100100;
		b = 32'b10100100010000001101101101001111;
		correct = 32'b00000100010000000001100001000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011010101011111001011100010;
		b = 32'b10001101000111110111110010111001;
		correct = 32'b00000001000101010111000010100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101111001111011110010100010;
		b = 32'b10000110101000010001010001110111;
		correct = 32'b00000100101000010001010000100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101001010000101001110111011;
		b = 32'b01010001111001111100101011110011;
		correct = 32'b00010001001000000100001010110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101110011001011011000010111;
		b = 32'b01101111010011100110110000000101;
		correct = 32'b00001101010011000010010000000101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100100010011011100011111110;
		b = 32'b10100011101000111000111111111001;
		correct = 32'b10000000100000011000100011111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111110100000100111100010011;
		b = 32'b11100010011100001111101010011001;
		correct = 32'b00000010010100000100101000010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111100101011010101111100011;
		b = 32'b01001111110011101110101110000000;
		correct = 32'b01000111100001001010101110000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010110100011101011010011010;
		b = 32'b01001110000100101011011000111011;
		correct = 32'b00001010000100001001011000011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111100110011010001010100000;
		b = 32'b00111010110110010110100001100011;
		correct = 32'b00001010100110010010000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000111000100000111100011100000;
		b = 32'b11110000011010001000000001110000;
		correct = 32'b10000000000000000000000001100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000000101010111101011001011;
		b = 32'b01010100101000100110010100000110;
		correct = 32'b00000000000000000110000000000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011100101011100011110100001;
		b = 32'b10100100010100010000010000000100;
		correct = 32'b10100000000100010000010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111100100101101011010010101;
		b = 32'b01110101000000101111110010001000;
		correct = 32'b00100101000000101101010010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000001101001010001001100001;
		b = 32'b10010111001010111111010001001110;
		correct = 32'b00000000001000001010000001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101001111100011111001110100;
		b = 32'b00110111000100001010111111011101;
		correct = 32'b00110101000100000010111001010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010110110001101111000111010;
		b = 32'b00000011110110101011000000011110;
		correct = 32'b00000010110110001001000000011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111100000011101110100000001;
		b = 32'b11111001111101101111001000001110;
		correct = 32'b00011001100000001101000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000001001000111110000010110;
		b = 32'b01000100111010011001010101001110;
		correct = 32'b00000000001000000001010000000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101011010010000100110001010;
		b = 32'b00101100011001011011011110001111;
		correct = 32'b00001100011000010000000110001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100000000110000111011110011;
		b = 32'b00100110111110000000001110101011;
		correct = 32'b00100100000000000000001010100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010101111111101100011111010;
		b = 32'b11110101011100001010101010101011;
		correct = 32'b11000000001100001000100010101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010010010010000111001101001;
		b = 32'b10100011100000000101000010001110;
		correct = 32'b00100010000000000000000000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111001100111100001111110110;
		b = 32'b00110100011001001010100111001011;
		correct = 32'b00100100001000001000000111000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111010100001010110001110110;
		b = 32'b10111111011101000010110000011110;
		correct = 32'b00100111010100000010110000010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000100000100010100100101101;
		b = 32'b10010010011111001111010001101111;
		correct = 32'b00000000000000000010000000101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101011000011100110001011000;
		b = 32'b10001010110011011001101000100110;
		correct = 32'b10001000010000011000100000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011110111100011011101011111;
		b = 32'b01101111111010111110110101011101;
		correct = 32'b01101011110010100010010101011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011011100100110111111000011;
		b = 32'b11000111100110001100001101101001;
		correct = 32'b00000011000100000100001101000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100001110100100001000001010;
		b = 32'b00100011110010011001100010000001;
		correct = 32'b00000000000010000000000000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001000000100100011111001001;
		b = 32'b01001010101011001001110100100111;
		correct = 32'b00001000000000000000010100000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101101101100001010100111001;
		b = 32'b11101101001101010011110001110111;
		correct = 32'b10000101001101000001010000110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000000011001011110110000000;
		b = 32'b00001111110001100110111100001110;
		correct = 32'b00001000000001000010110100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000101010110010111010010010;
		b = 32'b11010110010000100001010101110011;
		correct = 32'b00000000000000100000010000010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100101011000110010111110100;
		b = 32'b01011000101110000111100111000100;
		correct = 32'b00010000101010000110000111000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101000000000010001110101111;
		b = 32'b11000011010010111110011111000001;
		correct = 32'b00000001000000000010001110000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000011100100111111101000011;
		b = 32'b00010000011011110000000101011110;
		correct = 32'b00000000011000100000000101000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100010100110000000001010100;
		b = 32'b00000011100010001000100100011001;
		correct = 32'b00000000000000000000000000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011110100110101001011000010;
		b = 32'b01011111100001101001111010010111;
		correct = 32'b01010011100000100001001010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110110011101001001100111010;
		b = 32'b00011001100110011111110010101111;
		correct = 32'b00011000100010001001000000101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011111110100100110001110111;
		b = 32'b11110101110101101101100001100000;
		correct = 32'b11100001110100100100100001100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111000001010110010010000011;
		b = 32'b00101000011011110000110001011111;
		correct = 32'b00000000000001010000010000000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010001110100011001010001110;
		b = 32'b01011101001011000010110010011010;
		correct = 32'b01001000001010000010000010001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000000101000000101111010000;
		b = 32'b11011011100001000000110011001110;
		correct = 32'b01001000000001000000100011000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111010010011001010101010111;
		b = 32'b10101101111101001101100000000110;
		correct = 32'b00100101010000001001000000000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001110011101011100101010000;
		b = 32'b10010001111000110100100111111101;
		correct = 32'b00000001110000100000100101010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011011001010100101100111101;
		b = 32'b00010110001101111001100111111101;
		correct = 32'b00010010001001010000100100111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111011100000100110001010000;
		b = 32'b11000101000001001000101001000101;
		correct = 32'b11000101000000000000100001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011001110101010101000010110;
		b = 32'b00000101110101001010110010110111;
		correct = 32'b00000001000100001010100000010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000101101001000100100010111;
		b = 32'b11001101100101001010100110001011;
		correct = 32'b10000000100101001000100100000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010010000010011001000100101;
		b = 32'b11001101101000010011101010011000;
		correct = 32'b10001000000000010011001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111000100101110000010101100100;
		b = 32'b11010001010100001000101100111010;
		correct = 32'b00010000000100000000000100100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110111110000001101100010111;
		b = 32'b11010111110110000011101101001011;
		correct = 32'b01010110110110000001101100000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000000111011011011101010110;
		b = 32'b01100000001101010010110100000000;
		correct = 32'b01100000000101010010010100000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110111111011100110110111010;
		b = 32'b10110110000010001111010111001000;
		correct = 32'b10000110000010001100010110001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100100111100011010010110100;
		b = 32'b10000100001000011001111111001101;
		correct = 32'b10000100000000000001010010000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100001111100000111000010000;
		b = 32'b10000000100100100110011000110011;
		correct = 32'b10000000000100100000011000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011110010100000111000101100;
		b = 32'b11110111001111001011110010001010;
		correct = 32'b00010011000010000000110000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010000101101001111100111101;
		b = 32'b11001011111110011001110101101011;
		correct = 32'b10000010000100001001110100101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111110001000111100010001110;
		b = 32'b11111010111100000011100110110111;
		correct = 32'b01100010110000000011100010000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011000101001100010011001001;
		b = 32'b00100111001001000001100001101010;
		correct = 32'b00000011000001000000000001001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010010011111100001010000101;
		b = 32'b00010100010010010010111010100010;
		correct = 32'b00000000010010010000001010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000011111010001010001111111;
		b = 32'b01100010111111110000000001001110;
		correct = 32'b00100000011111010000000001001110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000010110001100000100010101111;
		b = 32'b01111001100100111010100111001110;
		correct = 32'b00000000100000100000100010001110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011111000110000010110000011;
		b = 32'b10000011001010101100000101000010;
		correct = 32'b00000011001000100000000100000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000000110110100100001011000;
		b = 32'b01010000000111000100101011110111;
		correct = 32'b00010000000110000100100001010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011011111110001000010000011;
		b = 32'b01100111101010101011111010100010;
		correct = 32'b00000011001010100001000010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011100101100011001010000000;
		b = 32'b00011001001110011111001001110000;
		correct = 32'b00010001000100000011001000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100110010110000010011111111;
		b = 32'b01110010001010001101000100001001;
		correct = 32'b01100000000010000000000000001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010110011000101001001100101;
		b = 32'b00100100111000111100110001101101;
		correct = 32'b00000000110000000100000001100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100100000010000010111010100;
		b = 32'b11011001110100000111101101000101;
		correct = 32'b11010000100000000000000101000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001110111001100000010111000;
		b = 32'b10110111000001011010000110011010;
		correct = 32'b00000001000001001000000010011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100101110111010101101110011;
		b = 32'b11100000101111101101000100110101;
		correct = 32'b11000000101110101000000100110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000101100111011000011010000;
		b = 32'b10010010111010011001010110111111;
		correct = 32'b10000000101000011001000010010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001111100010110101111011011;
		b = 32'b10010100110110011111110000110001;
		correct = 32'b00010000110100010110100000010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100101100111011000010111110;
		b = 32'b10111011110001110000100101001011;
		correct = 32'b00010000100000110000000000001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010000101110110011001101101;
		b = 32'b01100011110101010001011111111011;
		correct = 32'b00000010000101010000011001101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001010110100010111000111001;
		b = 32'b01111100111110011110111101111000;
		correct = 32'b01101000010110000010111000111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011000110010001010000100011;
		b = 32'b01011110010010100010010110001101;
		correct = 32'b00011010000010000000010000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000111010000100111001110010;
		b = 32'b11000011010000010100010000010100;
		correct = 32'b10000000010000000100010000010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001010011000000010110000001;
		b = 32'b10001111111000000110010001101110;
		correct = 32'b00000001010000000000010000000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110000111101111000001101001;
		b = 32'b11010011010111000011111000100000;
		correct = 32'b00010010000111000011000000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100001100111011100010011100;
		b = 32'b00110101011111111011101011100100;
		correct = 32'b00110100001100111011100010000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000000001111100101101011011;
		b = 32'b01001000001111001100000101011110;
		correct = 32'b00000000000001001100000101011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001110100111011110001111101;
		b = 32'b00101111101101100110010001100100;
		correct = 32'b00100001100100100010010001100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100011001011010010001111000;
		b = 32'b00100010101001000101000101101101;
		correct = 32'b00100000001001000000000001101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001011011101001000001011001;
		b = 32'b10010110010100100000111110111101;
		correct = 32'b00000000010000100000000000011001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111010010011001010111010111;
		b = 32'b01101101010100010110110100100111;
		correct = 32'b00101101010000010000010100000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101000000001001110101000100;
		b = 32'b10001100011011110010000101001101;
		correct = 32'b10000100000000000000000101000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000111100110100111000110001;
		b = 32'b01101101001101101110001100001111;
		correct = 32'b00000000001100100100001000000001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110011110010001011001001000;
		b = 32'b01000111010110010001011101110100;
		correct = 32'b00000110010110010001011001000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111011101000110010000111010;
		b = 32'b11011100000010011011110100110001;
		correct = 32'b00001100000000000010010000110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110000100110110011010011111;
		b = 32'b00100010000111001000111000101100;
		correct = 32'b00000010000100000000011000001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011110010100100011111101100;
		b = 32'b01111111110111110011001111000001;
		correct = 32'b01110011110010100000001111000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010111001011000100010010101;
		b = 32'b00000011000110000011001011101010;
		correct = 32'b00000010000000000000000010000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101011011000010100011010110;
		b = 32'b11010101001001000101101101000111;
		correct = 32'b00000101001001000000100001000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001111000011111001101011011;
		b = 32'b11001011110011111001011010001010;
		correct = 32'b00000001110000011001001000001010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110001110110011101011110110;
		b = 32'b10110000111000111001011011011101;
		correct = 32'b00010000001000110001001011010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100110100110001000100001110;
		b = 32'b00111100010010011010001011001000;
		correct = 32'b00011100010000010000000000001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001101000111001000010111000000;
		b = 32'b10001110110101000110111101000011;
		correct = 32'b00001100000101000000010101000000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101011011010010001110111000;
		b = 32'b11100011011010000101100110100011;
		correct = 32'b01000001011010000000000110100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011001010101010001110010010;
		b = 32'b01100001110001111101101010010001;
		correct = 32'b00100001000000101000001010010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001000110110101011111001000;
		b = 32'b11001110011111101011010100101010;
		correct = 32'b01000000000110100001010100001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000111000101000000110100011;
		b = 32'b10011100010000011100010010100111;
		correct = 32'b10000000010000001000000010100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001101100110110010110010100;
		b = 32'b01001011110111010011100101111111;
		correct = 32'b01001001100100010010000100010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101100100101100110011101100;
		b = 32'b00011001000111010000010000100001;
		correct = 32'b00000001000100000000010000100000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110100100000101011111111100;
		b = 32'b11000001111011111000000101101001;
		correct = 32'b01000000100000000000000101101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end

endmodule
