
    `include "alu.v"


    module mul_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .A(a),
                .B(b),
                .OpCode(op),
                .O(out)
            );
        /* create a 10Mhz clock */
        always
        #100 clock = ~clock; // every 100 nanoseconds invert
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, a, b, op, out);
            clock = 0;

    op = 3'b011;

		/* Display the operation */
		$display ("Opcode: 011, Operation: MUL");
		/* Test Cases!*/
		a = 32'b00001001111010001000001111111101;
		b = 32'b01101111100001111011001011000110;
		correct = 32'b00111001111101100111111111110100;
		#400 //5.597609e-33 * 8.39932e+28 = 0.0004701611
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110011010110001111101001100;
		b = 32'b11000100100010001000010100100000;
		correct = 32'b01100011011110101100010111001010;
		#400 //-4.235586e+18 * -1092.1602 = 4.6259382e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110011010000110000001010100;
		b = 32'b11010010111000010100010010100110;
		correct = 32'b10011001110011000111101011111010;
		#400 //4.370512e-35 * -483759700000.0 = -2.1142775e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111111011110010111100110000;
		b = 32'b01110000000000100101001100001010;
		correct = 32'b11111111111011110010111100110000;
		#400 //nan * 1.6133376e+29 = nan
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101101010000011100101111011100;
		b = 32'b10111100000001010001010001111001;
		correct = 32'b10101001110010010111110011010010;
		#400 //1.1016046e-11 * -0.008122557 = -8.947846e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000010111101111001110010100;
		b = 32'b11001101111111100011101001101011;
		correct = 32'b11111110110111010110100010001101;
		#400 //2.7600056e+29 * -533155170.0 = -1.4715112e+38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110111000111100010011000010;
		b = 32'b11100111001110010001001110111111;
		correct = 32'b01100110101001001010101011000010;
		#400 //-0.44486052 * -8.7400205e+23 = 3.88809e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010010011010010111111010101;
		b = 32'b11110100101100111011011111011000;
		correct = 32'b01011111100100000000101111001100;
		#400 //-1.8224253e-13 * -1.139099e+32 = 2.0759228e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101111001010110111100010100;
		b = 32'b11010011101111100101011111001110;
		correct = 32'b10101010001010101001011100100010;
		#400 //9.2667614e-26 * -1635033800000.0 = -1.5151468e-13
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110111100111101000111111001;
		b = 32'b11110011011111100011011110011101;
		correct = 32'b01111010111100100001111101001101;
		#400 //-31208.986 * -2.0141165e+31 = 6.2858535e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010000101111011100011111011;
		b = 32'b00111011110101001111010110111110;
		correct = 32'b10000110011111000110110110101001;
		#400 //-7.3051765e-33 * 0.0064990213 = -4.7476498e-35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001001011000101001011111000;
		b = 32'b00010010001010001011111010100011;
		correct = 32'b10111011111000110010110110001100;
		#400 //-1.3020441e+25 * 5.324643e-28 = -0.00693292
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101101001001111110000111010;
		b = 32'b01000100011110111101111011100000;
		correct = 32'b01101010101000100101001011110000;
		#400 //9.739011e+22 * 1007.4824 = 9.811882e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000011001000101100111101010;
		b = 32'b11000000101101101001010100111001;
		correct = 32'b00101001101000101101110100001000;
		#400 //-1.26760395e-14 * -5.7057157 = 7.232588e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111011001100010101101000000;
		b = 32'b11100100100001101110000001111100;
		correct = 32'b10111100011100101000100011110010;
		#400 //7.4371597e-25 * -1.9904316e+22 = -0.014803158
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100110010001100110000110010;
		b = 32'b10100011000010100011110000110000;
		correct = 32'b11100000010110001101101010010001;
		#400 //8.3408076e+36 * -7.49374e-18 = -6.2503845e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111010111011100010001100110;
		b = 32'b11011000011010110000110011111010;
		correct = 32'b11110000010010111001111010000111;
		#400 //243835600000000.0 * -1033763870000000.0 = -2.5206842e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000101011011111010001110111;
		b = 32'b01001101001011100101000011010001;
		correct = 32'b10100110011011001110011000100111;
		#400 //-4.49663e-24 * 182783250.0 = -8.2190863e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101011101110011011001101110;
		b = 32'b01000110010011111000011110101111;
		correct = 32'b01101100010010000110100000001010;
		#400 //7.2964286e+22 * 13281.921 = 9.691059e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001011010010010001011000000;
		b = 32'b01000000000100011000011110111110;
		correct = 32'b00010010000001001000100001001101;
		#400 //1.8391167e-28 * 2.27391 = 4.181986e-28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001110111000110011100010000;
		b = 32'b01000010011101111010001110111110;
		correct = 32'b10111100110101010011010001101010;
		#400 //-0.00042038457 * 61.909904 = -0.02602597
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000100010011111011000111101;
		b = 32'b00101101011100010100110000001001;
		correct = 32'b00011110100000100000100111001001;
		#400 //1.0038047e-09 * 1.3716147e-11 = 1.3768332e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010111010111000000100011011;
		b = 32'b00110101001110000001000101100001;
		correct = 32'b00010000101010010101010011001000;
		#400 //9.74023e-23 * 6.857063e-07 = 6.678937e-29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000100011100011100111000111110;
		b = 32'b11101000111100000011101001100110;
		correct = 32'b00101101111000101110100010000011;
		#400 //-2.8424116e-36 * -9.075562e+24 = 2.5796481e-11
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000010111001111100100001010;
		b = 32'b10100101010000110000110110001100;
		correct = 32'b00010110001010000101110101100100;
		#400 //-8.038944e-10 * -1.6918144e-16 = 1.3600401e-25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000111001010010100101011010;
		b = 32'b10000101000101111000010001110101;
		correct = 32'b10010110100001111010000111110110;
		#400 //30757540000.0 * -7.1243144e-36 = -2.1912638e-25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100101011010011010100011001;
		b = 32'b00101000100111011010010000000011;
		correct = 32'b10010101110101010101000100010001;
		#400 //-4.9228508e-12 * 1.750163e-14 = -8.6157915e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101110011001010110100101110;
		b = 32'b00111010110000011111101100111001;
		correct = 32'b00000001000110110001011101101011;
		#400 //1.9247684e-35 * 0.0014799602 = 2.8485805e-38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011101001101001110010100010;
		b = 32'b01001101111010001010111111100101;
		correct = 32'b01101010000101110111000001101101;
		#400 //9.379413e+16 * 487980200.0 = 4.576968e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110001011000000111000111101;
		b = 32'b01100000100011010001010110000011;
		correct = 32'b11100111001111011010010010011010;
		#400 //-11011.56 * 8.132941e+19 = -8.955636e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010000000001110100010011011;
		b = 32'b10100011100101110001101111110100;
		correct = 32'b11010110000110000010111010001110;
		#400 //2.5532982e+30 * -1.6383291e-17 = -41831430000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110011010100101000111100011;
		b = 32'b00101111110000010101101100110101;
		correct = 32'b10110110101100001111101100111000;
		#400 //-14996.472 * 3.5171302e-10 = -5.2744545e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011100111110101011000110001;
		b = 32'b01001010111001111100000011011011;
		correct = 32'b10100111000100000011111011001111;
		#400 //-2.6360043e-22 * 7594093.5 = -2.0018063e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111111011000111100010001111;
		b = 32'b11110110011011001100111101101011;
		correct = 32'b01011110110110101011111010111100;
		#400 //-6.563387e-15 * -1.2007705e+33 = 7.881121e+18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011001000110111010111000101;
		b = 32'b01100011000010100001100001101010;
		correct = 32'b11110110101100000101101000100110;
		#400 //-702055500000.0 * 2.54741e+21 = -1.7884232e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100100100111011000101101100;
		b = 32'b01111101000000110101000010000101;
		correct = 32'b11010010000101111000010001111101;
		#400 //-1.4913187e-26 * 1.0909184e+37 = -162690710000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110000110111111011100111000;
		b = 32'b11110100110111001111101010101001;
		correct = 32'b01011011100001101010000100101011;
		#400 //-5.411147e-16 * -1.4006217e+32 = 7.578971e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001010001011011111111111111;
		b = 32'b00100000000000110101001000101101;
		correct = 32'b00000001110010101110000101110011;
		#400 //6.70003e-19 * 1.1123321e-19 = 7.4526585e-38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100000001010101010100000111;
		b = 32'b10111010110000010111111111010001;
		correct = 32'b00110111010010011000111101011001;
		#400 //-0.008137948 * -0.0014762824 = 1.2013909e-05
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110000001111111111111110100;
		b = 32'b11000101011111101011110100010111;
		correct = 32'b01101100000001110101010001101000;
		#400 //-1.6056024e+23 * -4075.818 = 6.544143e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000001110110010111111000100;
		b = 32'b10101100001010111001101100110010;
		correct = 32'b10110100111110101111010011000101;
		#400 //191679.06 * -2.4386712e-12 = -4.6744222e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111100011011011001111010001;
		b = 32'b11000110101010110001001100100100;
		correct = 32'b10101110101111010110001101101010;
		#400 //3.933032e-15 * -21897.57 = -8.6123844e-11
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010010000110111011001110100;
		b = 32'b01011000110010010011010011101110;
		correct = 32'b11100011100110011010000001101011;
		#400 //-3202461.0 * 1769833300000000.0 = -5.6678224e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101000010000100011000110110;
		b = 32'b10111101100110011000111100010100;
		correct = 32'b11110011001000110111110001000000;
		#400 //1.7274815e+32 * -0.07497993 = -1.2952644e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001111100000011101001111011;
		b = 32'b00111101110101010001111000111110;
		correct = 32'b00001000010001111111110100001001;
		#400 //5.7832893e-33 * 0.10406159 = 6.0181826e-34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110110101010111100110011001;
		b = 32'b00100000000100001001110101110011;
		correct = 32'b01011111011100010010111101100011;
		#400 //1.4187847e+38 * 1.224937e-19 = 1.7379218e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111000110111100101011100101;
		b = 32'b01001100010110111001010001011111;
		correct = 32'b01111100000001011010000011011101;
		#400 //4.821546e+28 * 57561468.0 = 2.7753527e+36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110001011101010110000100011;
		b = 32'b00000100111101110110100111010001;
		correct = 32'b10111011101010001101000001001001;
		#400 //-8.856943e+32 * 5.8166598e-36 = -0.0051517827
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100010101011110111011111010;
		b = 32'b01111101010000000000001011100011;
		correct = 32'b01001010001000000111010110100101;
		#400 //1.6480838e-31 * 1.5951673e+37 = 2628969.2
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010110100111111101110000111;
		b = 32'b11111010111111110011100000111110;
		correct = 32'b01000110010100110101011000011110;
		#400 //-2.0413175e-32 * -6.625882e+35 = 13525.529
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011000010110111110001101001;
		b = 32'b11111010111001011000010010101001;
		correct = 32'b11010110011110100001110100100100;
		#400 //1.153801e-22 * -5.9586332e+35 = -68750766000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001011110011001110001011100;
		b = 32'b11101110101000000011111100000000;
		correct = 32'b01000000100111000011111100100111;
		#400 //-1.9690818e-28 * -2.4796882e+28 = 4.882709
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111000000001011101101101110;
		b = 32'b10000001100000100010110111101011;
		correct = 32'b10100001000000101110110010001010;
		#400 //9.276129e+18 * -4.7820347e-38 = -4.435877e-19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010100010001000100001100001;
		b = 32'b10110001111010110111000101010110;
		correct = 32'b11011100111110110010001101000110;
		#400 //8.252897e+25 * -6.852285e-09 = -5.6551202e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101110101000101100110111001;
		b = 32'b01001110011111100011001011111101;
		correct = 32'b11010100110100101101101101010001;
		#400 //-6795.2153 * 1066188600.0 = -7244981000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101110001000111100111011111;
		b = 32'b01000000101010101010100111111011;
		correct = 32'b11001111000000101111101101100011;
		#400 //-412040160.0 * 5.3332496 = -2197513000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000111111010000010000011001100;
		b = 32'b01010010011011010101111001000000;
		correct = 32'b10011010110101110011101111010011;
		#400 //-3.4926757e-34 * 254872130000.0 = -8.901857e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001100100101101110111100101;
		b = 32'b01110010011100111101001010010100;
		correct = 32'b01011100100010111110000101101111;
		#400 //6.522195e-14 * 4.8294036e+30 = 3.149831e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011100010000001110101110101;
		b = 32'b11000001000001001010001101011101;
		correct = 32'b01110101000011010000110000011001;
		#400 //-2.1568293e+31 * -8.289884 = 1.7879864e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011000000101001101011101010;
		b = 32'b01101000100010010001000111010000;
		correct = 32'b11110100000010111101101111111011;
		#400 //-8559338.0 * 5.1783423e+24 = -4.432318e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001011100011011010111001001;
		b = 32'b01101010110010010011010011000001;
		correct = 32'b01010100101111011111100110001010;
		#400 //5.3670423e-14 * 1.2162161e+26 = 6527483000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110000010001111001101010110;
		b = 32'b01100101011110101010010000100010;
		correct = 32'b10111100000001100001010101110000;
		#400 //-1.1062776e-25 * 7.397621e+22 = -0.008183822
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000011001010000100111010100;
		b = 32'b00111000100100011011101000000010;
		correct = 32'b11101001100000100110000011111100;
		#400 //-2.835358e+29 * 6.9487854e-05 = -1.9702294e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110101010001010001100111111;
		b = 32'b11010110111001101010100001110010;
		correct = 32'b10111110000101111111000110100001;
		#400 //1.170159e-15 * -126805570000000.0 = -0.14838268
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110111000001110101010000110;
		b = 32'b01111001110110000100100001100110;
		correct = 32'b01000001001111100000010101111101;
		#400 //8.4604036e-35 * 1.4037557e+35 = 11.87634
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011011100001111110001101011;
		b = 32'b11101110111010110101010101111100;
		correct = 32'b01010010110111011000100000101111;
		#400 //-1.3063878e-17 * -3.641616e+28 = 475736280000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101000101110001100011101111;
		b = 32'b01111011110110110110000000100000;
		correct = 32'b11111001100000010111101100010001;
		#400 //-0.036889013 * 2.2781253e+36 = -8.40378e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100001100111010000111110111;
		b = 32'b10011000101101110110110011111010;
		correct = 32'b00010101100000001011010100111111;
		#400 //-0.010963908 * -4.741443e-24 = 5.1984744e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010011110001001010101011110;
		b = 32'b01100101011000001011110001101010;
		correct = 32'b01001000010110100011100110100111;
		#400 //3.3689342e-18 * 6.6330357e+22 = 223462.61
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010001101111110000100111001;
		b = 32'b00011000001001000010011010010111;
		correct = 32'b00111010111010111101000000000001;
		#400 //8.479958e+20 * 2.1215986e-24 = 0.0017991067
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101111010001010011011010011;
		b = 32'b10101101000111101111110100101101;
		correct = 32'b11101011100100000111110100001100;
		#400 //3.8655887e+37 * -9.0374765e-12 = -3.4935167e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010100001101000011000110000;
		b = 32'b10010111010011110111001001000101;
		correct = 32'b11001010010110100000010100011010;
		#400 //5.3290514e+30 * -6.7029536e-25 = -3572038.5
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000010111010100000001100111;
		b = 32'b10100110110100001000000001110110;
		correct = 32'b11000111101101000011001101011010;
		#400 //6.3771424e+19 * -1.4467719e-15 = -92262.7
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011101110110010001010110110;
		b = 32'b11010001010111010101111100111011;
		correct = 32'b10110101101000011101001010010100;
		#400 //2.0289281e-17 * -59424092000.0 = -1.2056721e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011110001101100111011001011;
		b = 32'b00100110011000110110100101110100;
		correct = 32'b11010010101100001001101101000011;
		#400 //-4.8068773e+26 * 7.889936e-16 = -379259550000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101010010100001110111100011;
		b = 32'b11101010111110101001000100101000;
		correct = 32'b01111000110001011101001111001010;
		#400 //-211934770.0 * -1.5145847e+26 = 3.2099315e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001101010111100000100001111;
		b = 32'b00100101111011001000100001100111;
		correct = 32'b01100000000111101011000101111101;
		#400 //1.1147481e+35 * 4.1031904e-16 = 4.5740233e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010100100110101111101100011;
		b = 32'b00010010011110011010110010101111;
		correct = 32'b00111101100011111011101100110000;
		#400 //8.908127e+25 * 7.8783395e-28 = 0.07018125
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111101011101011110101110101;
		b = 32'b00010101001000110110010001100001;
		correct = 32'b00011101010111110000111001001011;
		#400 //89466.914 * 3.2996773e-26 = 2.9521194e-21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011011000101010110010010001;
		b = 32'b11010110100111000000101001001011;
		correct = 32'b01111010100010100010101001000110;
		#400 //-4.181399e+21 * -85784010000000.0 = 3.586972e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001001100001111110000001100;
		b = 32'b11110111100101011001010100001101;
		correct = 32'b01001001010011101101001101111101;
		#400 //-1.396162e-28 * -6.067776e+33 = 847159.8
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101110100011001010001111111;
		b = 32'b00111100011001111100110101000001;
		correct = 32'b00000010101111011100010100001000;
		#400 //1.9708814e-35 * 0.014148057 = 2.7884144e-37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001011111010100011000000100;
		b = 32'b10011011010000111010100010101010;
		correct = 32'b01010101010000011001001100110011;
		#400 //-8.219195e+34 * -1.618452e-22 = 13302372000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010011000010000010100011100;
		b = 32'b10000110100110000101101110100000;
		correct = 32'b10001001100001011110101110010010;
		#400 //56.25499 * -5.7310676e-35 = -3.2240115e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100100001011100110111111110;
		b = 32'b01001000010000100010110100011110;
		correct = 32'b01111101010010101111101101011111;
		#400 //8.480878e+31 * 198836.47 = 1.6863078e+37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000000101010101010100001010;
		b = 32'b11000111010000110110111110100100;
		correct = 32'b10100111111001000000000111001100;
		#400 //1.2648928e-19 * -50031.64 = -6.328466e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001101111011111101110111011;
		b = 32'b00001110111101001011110100011000;
		correct = 32'b00001001001101011010000001000011;
		#400 //0.00036236443 * 6.0332735e-30 = 2.1862437e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010011100100001011000010101;
		b = 32'b01110101110110110000110010000111;
		correct = 32'b11111000110011110010010010111101;
		#400 //-60.521564 * 5.5535503e+32 = -3.3610956e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101101100100000010111110110011;
		b = 32'b00100111001111111010111101111011;
		correct = 32'b00010101010101111110110011011001;
		#400 //1.6392087e-11 * 2.6601703e-15 = 4.3605744e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111110111011101100001011010;
		b = 32'b10101010100111001000000101011110;
		correct = 32'b00101011000001111001111111110010;
		#400 //-1.733165 * -2.7800933e-13 = 4.8183603e-13
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110101100000111101101010000;
		b = 32'b00010101111000101110001001101111;
		correct = 32'b00101101000111000110100011110110;
		#400 //97021835000000.0 * 9.163792e-26 = 8.890879e-12
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110011001010001010010001001;
		b = 32'b00111011011100100000110001101111;
		correct = 32'b11000010010110001001100010001010;
		#400 //-14661.134 * 0.003693368 = -54.148964
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100010101001010101001001101;
		b = 32'b10101001100000000000001110110101;
		correct = 32'b00001110010101001011000001110110;
		#400 //-4.6114422e-17 * -5.684985e-14 = 2.621598e-30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011010001100010100111100001;
		b = 32'b00111111010101101011000110110111;
		correct = 32'b10110011001001100011000010010011;
		#400 //-4.6138556e-08 * 0.8386492 = -3.8694065e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001100011010010100100100010;
		b = 32'b00110101111111100001011011111010;
		correct = 32'b01010000000011000001101101111011;
		#400 //4966649700000000.0 * 1.8931162e-06 = 9402445000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110100000101111010101110001;
		b = 32'b01111010001001110010100101111000;
		correct = 32'b01011001001010110000011010100111;
		#400 //1.3865798e-20 * 2.1698867e+35 = 3008721000000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111000111000010110101010111;
		b = 32'b00010001010010010100001010000011;
		correct = 32'b10101000111101011001000001011010;
		#400 //-171718550000000.0 * 1.58766e-28 = -2.7263067e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000000010101001110010000011;
		b = 32'b00001100000001110100011101011101;
		correct = 32'b00011100100100100111111001011010;
		#400 //9302052000.0 * 1.0421497e-31 = 9.694131e-22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011100001011001110010101101;
		b = 32'b10111000000110000010010001100001;
		correct = 32'b00110100000111101101000000000111;
		#400 //-0.004077515 * -3.6273505e-05 = 1.4790577e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100000010010010111100001111;
		b = 32'b10100010110010100101110101110100;
		correct = 32'b00110111010110001110001001101100;
		#400 //-2356800000000.0 * -5.4851157e-18 = 1.2927321e-05
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011010111001011100111101110;
		b = 32'b01100010101000110011011010000001;
		correct = 32'b10101110100011001011100101100001;
		#400 //-4.2510337e-32 * 1.5053734e+21 = -6.399393e-11
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111100011110010101001111110;
		b = 32'b01111101011101011100001010111000;
		correct = 32'b01110101100010010111000010010000;
		#400 //1.7066715e-05 * 2.0416994e+37 = 3.4845103e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101101100001001010011110100;
		b = 32'b01110110110101010011110101101010;
		correct = 32'b00111101000100110001011001001100;
		#400 //1.6605677e-35 * 2.1625095e+33 = 0.035909936
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011001100011101101011101110;
		b = 32'b00010001111001110010110000010111;
		correct = 32'b00110101101000001001101100101110;
		#400 //3.2808492e+21 * 3.6472546e-28 = 1.1966092e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110100011110000100110101000;
		b = 32'b01001011010100101000011010011110;
		correct = 32'b00110010011010110100001001000110;
		#400 //9.925236e-16 * 13797022.0 = 1.3693869e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011101100010010100010110001;
		b = 32'b01010101010110100011111111000100;
		correct = 32'b11110001100101110000100011000111;
		#400 //-9.973162e+16 * 14997963000000.0 = -1.4957711e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001110111110110111110100100;
		b = 32'b10100011011101110001111101100010;
		correct = 32'b00111101110101111011000000011011;
		#400 //-7861459000000000.0 * -1.3396542e-17 = 0.10531636
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100100110010000100011010000;
		b = 32'b11010100101111100011100111011101;
		correct = 32'b01111001111000110110111001000011;
		#400 //-2.2583895e+22 * -6536116600000.0 = 1.4761097e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000110101110010001011000111;
		b = 32'b00110100010000011101000101110000;
		correct = 32'b00001101101000101110000100111010;
		#400 //5.5611314e-24 * 1.8050719e-07 = 1.0038242e-30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000111000011110010101110011;
		b = 32'b01000000110000100000110110101000;
		correct = 32'b01010010001010110011101111101110;
		#400 //30319286000.0 * 6.064167 = 183861220000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101000111000001000111011010;
		b = 32'b11000011001011001001111011000000;
		correct = 32'b00101000110100100111100110001101;
		#400 //-1.3536891e-16 * -172.62012 = 2.3367398e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110111010100011101000010011;
		b = 32'b11011110001010000110011001011011;
		correct = 32'b10100101100110100001001111000011;
		#400 //8.810635e-35 * -3.0336216e+18 = -2.6728133e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010001011010001011010100110;
		b = 32'b10111111110010100001000101010100;
		correct = 32'b10000010100010001001111110010110;
		#400 //1.2716532e-37 * -1.5786538 = -2.0075002e-37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100011101000100100000101001;
		b = 32'b10100111001111010111011101010101;
		correct = 32'b11011100001101001100101100100101;
		#400 //7.7416017e+31 * -2.629371e-15 = -2.0355542e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011101111011110001110110010;
		b = 32'b11100010101100110100000011010110;
		correct = 32'b11111111000001001111011001001101;
		#400 //1.0689825e+17 * -1.6533196e+21 = -1.7673696e+38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111100001001001101100011000;
		b = 32'b00101100111001001101011110100001;
		correct = 32'b01010100111011010001001110100110;
		#400 //1.2524267e+24 * 6.5040894e-12 = 8145895000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000010111010110001111001111110;
		b = 32'b01000101110100110011111001110000;
		correct = 32'b10001001010000100000001101111010;
		#400 //-3.4547648e-37 * 6759.8047 = -2.3353535e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011101001110000000111000101;
		b = 32'b10101110100111111100011001110001;
		correct = 32'b10101010110100000111011100011101;
		#400 //0.0050966465 * -7.265733e-11 = -3.7030874e-13
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010101100010011100101101111;
		b = 32'b10101100010011101001001101100011;
		correct = 32'b10001111100011110000001001000000;
		#400 //4.8036756e-18 * -2.9356177e-12 = -1.4101755e-29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100001011101010111100001101;
		b = 32'b10001001111001100001110001101010;
		correct = 32'b00011110100111010000010010101001;
		#400 //-3001044700000.0 * -5.5397206e-33 = 1.6624949e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111101100001010011010100111;
		b = 32'b00000110001011001011101001111010;
		correct = 32'b10001110011011100110000101001011;
		#400 //-90445.305 * 3.2486606e-35 = -2.938261e-30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111011100100010101110010111;
		b = 32'b11111011101111010011010001001010;
		correct = 32'b11110011101100101111101110100101;
		#400 //1.4434473e-05 * -1.9648093e+36 = -2.8360986e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011100101010101101011011010;
		b = 32'b00111110001011011000000010011101;
		correct = 32'b11010010010010100111001011011101;
		#400 //-1282948700000.0 * 0.16943593 = -217377620000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000000000101011000010100010;
		b = 32'b00000000011010010100110001011000;
		correct = 32'b10010000110101110000010110101111;
		#400 //-8770456000.0 * 9.670114e-39 = -8.4811304e-29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001001001100000111101000100;
		b = 32'b10100000000001100110111110101010;
		correct = 32'b00100001101011100110100011011001;
		#400 //-10.378727 * -1.1387188e-19 = 1.1818452e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000101011010010000011100011;
		b = 32'b11111110100011001001111100011111;
		correct = 32'b11010111101111100011001100110001;
		#400 //4.475266e-24 * -9.345906e+37 = -418254150000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010000111011011000110001001;
		b = 32'b00110011011101111111001100001110;
		correct = 32'b10010110000110001011110000000011;
		#400 //-2.1371454e-18 * 5.7730226e-08 = -1.2337788e-25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100100010101000111011000111;
		b = 32'b11000010100000000110101101010010;
		correct = 32'b11110111100010110000001011110011;
		#400 //8.782139e+31 * -64.20961 = -5.638977e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000011100010110111110100111;
		b = 32'b10100011000111000011011010110010;
		correct = 32'b10000100000100110101001110011111;
		#400 //2.0450437e-19 * -8.468359e-18 = -1.7318164e-36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110010100111111101010101011;
		b = 32'b00001101100100000111001111000101;
		correct = 32'b10110100011011110011100110111010;
		#400 //-2.5026083e+23 * 8.902556e-31 = -2.227961e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010000111111001100010010011;
		b = 32'b11101001110111100100011101011110;
		correct = 32'b01011100100010101001001011001101;
		#400 //-9.2897094e-09 * -3.358982e+25 = 3.1203965e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000100110011001111000001110;
		b = 32'b11001110100001111000001000101101;
		correct = 32'b00101111101000101010000011101101;
		#400 //-2.60238e-19 * -1136727700.0 = 2.9581973e-10
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000100011101010100101011011;
		b = 32'b00000011001110111110111011111110;
		correct = 32'b00111100010100010111010111001001;
		#400 //2.314816e+34 * 5.522871e-37 = 0.01278443
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001000011010110110000000111;
		b = 32'b01110000101110000110101100001001;
		correct = 32'b11110010010010111100000110001100;
		#400 //-8.838874 * 4.565971e+29 = -4.0358042e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111001001010011100001110001;
		b = 32'b00010000011001111100101101110110;
		correct = 32'b11000000000101011001100100111110;
		#400 //-5.113326e+28 * 4.5713458e-29 = -2.3374782
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101000100011001111010110010;
		b = 32'b00101100100100011001000010011101;
		correct = 32'b01001010001001011001101001001011;
		#400 //6.5581374e+17 * 4.137203e-12 = 2713234.8
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001011110110001101110100011;
		b = 32'b01001010110000010000000110001111;
		correct = 32'b01000100101111010101000101011101;
		#400 //0.00023947521 * 6324423.5 = 1514.5426
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111000001110001111111110010;
		b = 32'b00110000001011101000001001111100;
		correct = 32'b00010111101110000011100100101100;
		#400 //1.8752331e-15 * 6.348626e-10 = 1.1905154e-24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000010101011010011110010001;
		b = 32'b00010001001010011111111011101001;
		correct = 32'b10100010000011011110000001011101;
		#400 //-14338115000.0 * 1.34103e-28 = -1.922784e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100110100011101001001111101;
		b = 32'b10111111100110100010101101111100;
		correct = 32'b01111100111111001011100010000110;
		#400 //-8.715674e+36 * -1.204452 = 1.0497611e+37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101000011001011000001101110;
		b = 32'b01110101101100110101010011110110;
		correct = 32'b11101011010001010001110000011100;
		#400 //-5.2410803e-07 * 4.5466033e+32 = -2.3829113e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000100111001101110000101000;
		b = 32'b11100101010010011111100100110100;
		correct = 32'b11100110011101111000001100011011;
		#400 //4.9018745 * -5.961204e+22 = -2.9221075e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011100001000001111011101001;
		b = 32'b11010011011010010101001011001100;
		correct = 32'b11000111011100001101010110111011;
		#400 //6.1523515e-08 * -1002116500000.0 = -61653.73
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011110010111101011110011111;
		b = 32'b00110001101101010111001110101010;
		correct = 32'b11000110000100000111101110001101;
		#400 //-1750991800000.0 * 5.280943e-09 = -9246.888
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110111110011011011101011100;
		b = 32'b00011001111101100100110011011001;
		correct = 32'b11010001011100000100000100101001;
		#400 //-2.5324236e+33 * 2.5466842e-23 = -64492835000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011111010010101010010110011;
		b = 32'b00110111111001000111111101000000;
		correct = 32'b01101100010100000100001101101011;
		#400 //3.697275e+31 * 2.7238973e-05 = 1.0070998e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000011010010110010011010011;
		b = 32'b10001110000101000000100000100101;
		correct = 32'b10110111000001101111010110110111;
		#400 //4.408685e+24 * -1.824633e-30 = -8.044232e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101010101111000111100000010;
		b = 32'b01000101010011111111101101100001;
		correct = 32'b11001011001011110010000001001110;
		#400 //-3448.938 * 3327.7112 = -11477070.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011011010000101000000001001;
		b = 32'b11101000111001110110111101110001;
		correct = 32'b01000100110100100000010101011001;
		#400 //-1.9216451e-22 * -8.743379e+24 = 1680.1671
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110110010000110000010001010;
		b = 32'b00010101111100111110110101110100;
		correct = 32'b10101101001111101110110101111111;
		#400 //-110158480000000.0 * 9.8521553e-26 = -1.0852984e-11
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000110110000011100011001010;
		b = 32'b01100011100001010101010100100001;
		correct = 32'b10110100111000010011101011001111;
		#400 //-8.5284475e-29 * 4.9191023e+21 = -4.1952305e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111010101110011011100110010111;
		b = 32'b10001110110000010111101011010011;
		correct = 32'b01001010000011000101111000000110;
		#400 //-4.8216956e+35 * -4.769645e-30 = 2299777.5
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011011011010100110110011011;
		b = 32'b01000100000001100011000101111111;
		correct = 32'b00101111111110001100100100000001;
		#400 //8.4307013e-13 * 536.7734 = 4.525376e-10
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011011100100001100111110010;
		b = 32'b10000010110101000011011011111100;
		correct = 32'b10011110110010001011000101111100;
		#400 //6.814547e+16 * -3.118216e-37 = -2.124923e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000100100100111101010101010;
		b = 32'b01000101010011100001001100101011;
		correct = 32'b01010110011010111101001101011001;
		#400 //19660100000.0 * 3297.198 = 64823240000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011100111011011000111101101;
		b = 32'b11000000101011111001001111100110;
		correct = 32'b10110100110110000100111101111000;
		#400 //7.343247e-08 * -5.486804 = -4.0290956e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100101010001000111010010101;
		b = 32'b01110100011111011001000110000000;
		correct = 32'b11110001101001101111010010110110;
		#400 //-0.0205758 * 8.035902e+31 = -1.6534512e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011100100011000100010011100;
		b = 32'b01001101011101100000101101111101;
		correct = 32'b01011001100010111101111111001110;
		#400 //19075384.0 * 257996750.0 = 4921387000000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010011100000100001000101001;
		b = 32'b01001010001011001100000010011000;
		correct = 32'b01010101001000100010000100110100;
		#400 //3936394.2 * 2830374.0 = 11141468000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100100100010111011110010100;
		b = 32'b00101101000010011010000101010010;
		correct = 32'b11100010000111000110100101010010;
		#400 //-9.220073e+31 * 7.823369e-12 = -7.213203e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100101011011010111001001111;
		b = 32'b01101110011101101111111000001011;
		correct = 32'b01100011101001111001000111011010;
		#400 //3.2350587e-07 * 1.9110108e+28 = 6.182232e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110111100011000000011000010;
		b = 32'b00011111110100001101101111111011;
		correct = 32'b10101111010001010000100000100100;
		#400 //-2025873700.0 * 8.8455354e-20 = -1.7919938e-10
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111110010100000100111100111;
		b = 32'b01001100110111011000111110011101;
		correct = 32'b11010101001011101101101111100100;
		#400 //-103443.805 * 116161770.0 = -12016215000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010011000010000001011011001;
		b = 32'b01100010000111110010100100000001;
		correct = 32'b10101101000010111110010011001111;
		#400 //-1.08338915e-32 * 7.3399674e+20 = -7.952041e-12
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110100000000111001111111010;
		b = 32'b00100010001000110100010011100100;
		correct = 32'b01010001001000111101100011010011;
		#400 //1.9877144e+28 * 2.212709e-18 = 43982336000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011111110010111101110000001;
		b = 32'b10100011111011100101100000011110;
		correct = 32'b00011000011010000100011010110010;
		#400 //-1.1617431e-07 * -2.584133e-17 = 3.002099e-24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010111000111001011011001110;
		b = 32'b10001000100100010110011011101100;
		correct = 32'b00110100000000010100001111101011;
		#400 //-1.3756916e+26 * -8.751067e-34 = 1.203877e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011101011000110010011001100;
		b = 32'b00100110110101000001110011110010;
		correct = 32'b11011011000011101101011011110111;
		#400 //-2.7316878e+31 * 1.4718301e-15 = -4.0205803e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011111011110010101110001110;
		b = 32'b11101110010001111101101101100001;
		correct = 32'b01111010101110101011011111010000;
		#400 //-31348508.0 * -1.5463182e+28 = 4.847477e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111001001101100101100011010;
		b = 32'b01011010111010100100000100011111;
		correct = 32'b10111010100110001010000000010100;
		#400 //-3.531987e-20 * 3.2968373e+16 = -0.0011644387
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011000000110000001100001110;
		b = 32'b01101101111100100100110000001100;
		correct = 32'b11100001011101111111111110011101;
		#400 //-3.0503593e-08 * 9.3734134e+27 = -2.859228e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100100110011110110000000000;
		b = 32'b11010010110101011101001001011010;
		correct = 32'b00101000000000001000111111010110;
		#400 //-1.5542138e-26 * -459178570000.0 = 7.136617e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111001000111110110111010101;
		b = 32'b00111110101001010110010011110011;
		correct = 32'b10011110010100111101000111011110;
		#400 //-3.4713323e-20 * 0.3230358 = -1.12136465e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110010101000110110110110101;
		b = 32'b00100010111000100110010111010110;
		correct = 32'b01000001101110111101110101011011;
		#400 //3.8267724e+18 * 6.1365246e-18 = 23.483084
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111101111100111001111101001;
		b = 32'b11001110100010111010000011111001;
		correct = 32'b00011110110011111100000101100010;
		#400 //-1.8780093e-29 * -1171291300.0 = 2.1996959e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010001001110011000011011011;
		b = 32'b10100001010000111000011001010101;
		correct = 32'b10111011111111110110001111100100;
		#400 //1.176501e+16 * -6.6246357e-19 = -0.0077938903
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011010000110100000100101001;
		b = 32'b10000011011011110111101100101101;
		correct = 32'b00111111001101101010011111001000;
		#400 //-1.0138195e+36 * -7.0377186e-37 = 0.71349764
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001000001101010101011111111;
		b = 32'b01000111011000001100100100101111;
		correct = 32'b10001000111011000111111011101000;
		#400 //-2.4734597e-38 * 57545.184 = -1.4233569e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010111100110100111110110110;
		b = 32'b00010100100101001111001001010111;
		correct = 32'b00100000000011011001000001101001;
		#400 //7972827.0 * 1.5039767e-26 = 1.1990946e-19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011110011101010010010110001;
		b = 32'b00111110111011101010010011010001;
		correct = 32'b11101011010000001010001000100111;
		#400 //-4.996329e+26 * 0.4661012 = -2.328795e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000000011100111011111011111;
		b = 32'b01000010101101011101100010110001;
		correct = 32'b10011011010010100110011010110001;
		#400 //-1.841359e-24 * 90.923225 = -1.674223e-22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100111111000000101011011101;
		b = 32'b01000100010100101001011001001011;
		correct = 32'b11001001110011110101010011100001;
		#400 //-2016.3395 * 842.3483 = -1698460.1
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001111011000110000001000000;
		b = 32'b10100000001000010011111010111110;
		correct = 32'b11000010100101001110001001110111;
		#400 //5.450459e+20 * -1.365799e-19 = -74.442314
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000011000000001110000110011;
		b = 32'b00011111100010000010101010010000;
		correct = 32'b11000000011011100110100001111100;
		#400 //-6.4595354e+19 * 5.7668654e-20 = -3.7251272
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011001000001101011100010101;
		b = 32'b01001000000101010111100000010110;
		correct = 32'b00010011101110111101000101000100;
		#400 //3.097669e-32 * 153056.34 = 4.741179e-27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001011101111001100100010000;
		b = 32'b10011101001110101010000010000100;
		correct = 32'b10001111001101001000000001110101;
		#400 //3.6030237e-09 * -2.469988e-21 = -8.899425e-30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100100001110101001111010001;
		b = 32'b11100011011110111011010000010111;
		correct = 32'b01111000100001010000111001100001;
		#400 //-4649814300000.0 * -4.6431096e+21 = 2.1589598e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010010101110010101111110101;
		b = 32'b11000001110100010100100111011111;
		correct = 32'b01011100101011111110100011111010;
		#400 //-1.5141363e+16 * -26.16107 = 3.9611425e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111111011101111110001011000;
		b = 32'b10001001110110100011101001001011;
		correct = 32'b10111010010010111011100101001110;
		#400 //1.4792499e+29 * -5.253641e-33 = -0.0007771448
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000001110100111011001101001;
		b = 32'b11000011000111000001100100110010;
		correct = 32'b00010011111000110110010100000100;
		#400 //-3.6773252e-29 * -156.09842 = 5.7402465e-27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000011101000001011011000001;
		b = 32'b01000000011111110000011111100100;
		correct = 32'b10011001011100110010101000110000;
		#400 //-3.1547749e-24 * 3.9848566 = -1.2571325e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001001010011001010010110001;
		b = 32'b11010010011100001100010000110010;
		correct = 32'b01000100000111110111110101011101;
		#400 //-2.4677258e-09 * -258520940000.0 = 637.9588
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110101101000100101111111101;
		b = 32'b10100011011100110101011101001000;
		correct = 32'b00111010101010110110000110011010;
		#400 //-99119230000000.0 * -1.3191539e-17 = 0.0013075352
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001001111001010110100101111;
		b = 32'b10100111100000011101001011001110;
		correct = 32'b11100001001111110101110101000101;
		#400 //6.1229024e+34 * -3.6033247e-15 = -2.2062806e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111001011011101001110110101;
		b = 32'b01011000001101101100111010010101;
		correct = 32'b11110111111110000100000110010000;
		#400 //-1.2525554e+19 * 803993500000000.0 = -1.0070464e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111101011001100101110100110;
		b = 32'b10011010011011110010001111111101;
		correct = 32'b10001010101000010110101001101011;
		#400 //3.143132e-10 * -4.9453113e-23 = -1.5543766e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000010001100000011001111001;
		b = 32'b00110100100101000001101111100100;
		correct = 32'b11011101011001010010001010100010;
		#400 //-3.7405919e+24 * 2.758744e-07 = -1.0319336e+18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001001101000001110111000001;
		b = 32'b10100110000111101100010010011001;
		correct = 32'b00100111110111110110100101011111;
		#400 //-11.257264 * -5.50837e-16 = 6.2009177e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111011000010011010010001101;
		b = 32'b11001100001110000010000110110100;
		correct = 32'b10011100001000011111101101101011;
		#400 //1.11034774e-29 * -48269010.0 = -5.359538e-22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101111001011100001111111100;
		b = 32'b00110110011100111011100011111010;
		correct = 32'b00110100110110101011111100001101;
		#400 //0.11219022 * 3.6317492e-06 = 4.0744672e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000010110010011001011100111;
		b = 32'b10111110000010011010011110000100;
		correct = 32'b00111110111010011001010010111100;
		#400 //-3.3937318 * -0.13442808 = 0.45621288
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010000101110100011000001010;
		b = 32'b11111011101000110000110001000100;
		correct = 32'b01001110010000001011000110110000;
		#400 //-4.773353e-28 * -1.6931863e+36 = 808217600.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100010110000110101000111001;
		b = 32'b10100101000000011010110000000011;
		correct = 32'b00001001110110110011110111100001;
		#400 //-4.6927508e-17 * -1.1247246e-16 = 5.2780523e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011101111100011010011110111;
		b = 32'b10111011110000000001010011100100;
		correct = 32'b00010000000011101011011100111111;
		#400 //-4.801497e-27 * -0.0058618654 = 2.814573e-29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010010001111110100100100010;
		b = 32'b00110100010000101101010100110010;
		correct = 32'b01011111000110000010010100101000;
		#400 //6.0419294e+25 * 1.8145218e-07 = 1.0963213e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100011000011111011010101101;
		b = 32'b01010100011001001000000000010000;
		correct = 32'b01110001010010011011000010111100;
		#400 //2.5441237e+17 * 3925604300000.0 = 9.987223e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000111101111011111000010010;
		b = 32'b10101010111011000110100011100000;
		correct = 32'b00011100011001001100100010110111;
		#400 //-1.8025637e-09 * -4.1994793e-13 = 7.569829e-22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111001110000010101000011001;
		b = 32'b10101110010001101010001110010000;
		correct = 32'b01000110000011101110011000111010;
		#400 //-202490950000000.0 * -4.516526e-11 = 9145.557
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000101011011101100000100011;
		b = 32'b10110101111000001001011101101000;
		correct = 32'b11001111000110001000001111110000;
		#400 //1529150500000000.0 * -1.6733366e-06 = -2558783500.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011110101110101011101100100;
		b = 32'b10101101110111101101001110110100;
		correct = 32'b01101010001110110110111111011101;
		#400 //-2.2362326e+36 * -2.5332493e-11 = 5.6649347e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101100011010000101010111111;
		b = 32'b11010111010010000011110010110001;
		correct = 32'b11011101010111001010001110101011;
		#400 //4513.3433 * -220163000000000.0 = -9.936712e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011000000000101111001000001;
		b = 32'b11001111110000000110101011000010;
		correct = 32'b10110011010000001111100001110010;
		#400 //6.958853e-18 * -6456444000.0 = -4.4929443e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001000111110010111000010111;
		b = 32'b00000110001110001101100101101101;
		correct = 32'b00111111111001011110000010100101;
		#400 //5.1656876e+34 * 3.4766293e-35 = 1.7959181
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101100111010111010101100110;
		b = 32'b10011100111100001010101111100111;
		correct = 32'b00100011000101000000011111001011;
		#400 //-5038.675 * -1.5926303e-21 = 8.024746e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010101011101000110011001001;
		b = 32'b00110111111000010111010101110110;
		correct = 32'b00111011000110011011100111010011;
		#400 //87.27497 * 2.6876787e-05 = 0.0023456707
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101101110100110110001110111;
		b = 32'b01100111101111101110110100111001;
		correct = 32'b00111110000010110000100101000000;
		#400 //7.529593e-26 * 1.8032512e+24 = 0.13577747
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110000101110001101001110001;
		b = 32'b00010100100100101110111111011010;
		correct = 32'b00011011001011010111010101001110;
		#400 //9670.61 * 1.4836837e-26 = 1.4348128e-22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100101100111000101000110001;
		b = 32'b01010010001100011111100011001100;
		correct = 32'b00010111011110011010001000010010;
		#400 //4.2209607e-36 * 191095830000.0 = 8.06608e-25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001000010001001001000011010;
		b = 32'b10010001011011000011001010001000;
		correct = 32'b00110010111111000000001101001010;
		#400 //-1.574553e+20 * -1.8632689e-28 = 2.9338157e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100110011000101010100111100;
		b = 32'b01011100110000010011111010000000;
		correct = 32'b01000010000110100011111000100101;
		#400 //8.861529e-17 * 4.3514712e+17 = 38.560688
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101101110000001101000101111;
		b = 32'b11010111000000101010110101010110;
		correct = 32'b00111101001110111111001111100111;
		#400 //-3.1936655e-16 * -143680980000000.0 = 0.0458869
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100011000001100001100011101;
		b = 32'b00101101000011001010110110000001;
		correct = 32'b00110001111101110000011000010010;
		#400 //899.04865 * 7.996604e-12 = 7.1893362e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111010000101000000110110111;
		b = 32'b00001010000010110100001111100011;
		correct = 32'b11000001110100111010000000000110;
		#400 //-3.9450645e+33 * 6.7053746e-33 = -26.453136
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101000000010001100010000101;
		b = 32'b11100100110111101011110001000000;
		correct = 32'b11001010011000001010010001100011;
		#400 //1.1197274e-16 * -3.2869936e+22 = -3680536.8
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110110010011010111010011000;
		b = 32'b11001011011101011110101010010010;
		correct = 32'b00011010110000011011110011100100;
		#400 //-4.9718453e-30 * -16116370.0 = 8.01281e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000001111011010010000001001;
		b = 32'b01110001000111011001101011011101;
		correct = 32'b11010001111010011000000010100100;
		#400 //-1.6063197e-19 * 7.804218e+29 = -125360700000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111111011111001000000101101;
		b = 32'b01000011110111100001111010100100;
		correct = 32'b00101100010011111101101110110011;
		#400 //6.649214e-15 * 444.23938 = 2.9538427e-12
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101111001000101010011111110;
		b = 32'b11110110110010000111001101100101;
		correct = 32'b11011101001100101100100101010011;
		#400 //3.9609288e-16 * -2.0328122e+33 = -8.051825e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101010000100010000001100001001;
		b = 32'b00100100010110010001011011001001;
		correct = 32'b11001110111101011111000011110101;
		#400 //-4.3827144e+25 * 4.7073674e-17 = -2063104600.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011101000010001001011011001;
		b = 32'b11010001000101110110110111000010;
		correct = 32'b11110101001111101000111001011010;
		#400 //5.942568e+21 * -40648843000.0 = -2.415585e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110111001010111111001100111111;
		b = 32'b00000010001010100001001001010001;
		correct = 32'b00111001111001000111011110101011;
		#400 //3.487564e+33 * 1.2494884e-37 = 0.00043576708
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001100001001111111111101100;
		b = 32'b01011001100111111110011100110111;
		correct = 32'b11111011101001100010011000100110;
		#400 //-3.066764e+20 * 5626093000000000.0 = -1.72539e+36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001000000100110000001001001;
		b = 32'b01001101110010011101111000010001;
		correct = 32'b01100111010011011001110101100011;
		#400 //2293600900000000.0 * 423346720.0 = 9.709884e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000101000110110100110000100;
		b = 32'b00101110100000110101100000010101;
		correct = 32'b01010111101001111010111001110000;
		#400 //6.173537e+24 * 5.972837e-11 = 368735300000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111000110000101011100011111;
		b = 32'b00111010101001110010101100100010;
		correct = 32'b00100010010001101111010100000000;
		#400 //2.1141466e-15 * 0.0012753943 = 2.6963706e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110111011111010100100000001011;
		b = 32'b10001000001001100001111001001001;
		correct = 32'b11000000001001000101101010101110;
		#400 //5.1371575e+33 * -4.998941e-34 = -2.5680346
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101100001111001011010001000;
		b = 32'b11000011111000110001001101111010;
		correct = 32'b00001001111100001000100110010111;
		#400 //-1.2750635e-35 * -454.15216 = 5.7907287e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010011011110101001110110100;
		b = 32'b11100101100011001001001000100110;
		correct = 32'b01011000100000110110101001101000;
		#400 //-1.3930663e-08 * -8.297841e+22 = 1155944300000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010110101110101100110000001;
		b = 32'b00110110001000101100110101000001;
		correct = 32'b00110001100010001111001101001101;
		#400 //0.0016429872 * 2.4259355e-06 = 3.985781e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000000110101011011110001000;
		b = 32'b11101101010001100001010011000100;
		correct = 32'b01011101111011110110110100000000;
		#400 //-5.6285687e-10 * -3.831446e+27 = 2.1565557e+18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110110001000101010111000001;
		b = 32'b01011011110011001111100000101001;
		correct = 32'b01010011000111010011001010101000;
		#400 //5.8512383e-06 * 1.153875e+17 = 675159740000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101101011101001000011001010;
		b = 32'b00111010001011010001111101011001;
		correct = 32'b01100000011011000001101001110001;
		#400 //1.0304533e+23 * 0.00066040974 = 6.805214e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100100101101001111111110000;
		b = 32'b00111001000110010000100100011010;
		correct = 32'b10001110001101000001010111100011;
		#400 //-1.5209214e-26 * 0.00014594608 = -2.2197251e-30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001101010001001111111101111;
		b = 32'b00110111101100101001110101100110;
		correct = 32'b00000001111010110100110111000011;
		#400 //4.059493e-33 * 2.1292548e-05 = 8.643695e-38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001011101110000111010010100;
		b = 32'b11110001111011101011010100000111;
		correct = 32'b01001011111001100101111001000010;
		#400 //-1.2772545e-23 * -2.364041e+30 = 30194820.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110100111011011110101011001;
		b = 32'b01111010011110000111000010101110;
		correct = 32'b11010001100110010001010011011100;
		#400 //-2.5484213e-25 * 3.2249376e+35 = -82184995000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101111011011011010101101101;
		b = 32'b11000100100111110011111101100111;
		correct = 32'b10001011000100111101111010001110;
		#400 //2.2354018e-35 * -1273.9813 = -2.8478602e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001001011101110111000110111;
		b = 32'b00001001001100110110111101011000;
		correct = 32'b00010010111101010011100101001100;
		#400 //716515.44 * 2.1598695e-33 = 1.54757985e-27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011111011000011001100010010;
		b = 32'b11000011110111110110110100100110;
		correct = 32'b00010000010011100010010100110001;
		#400 //-9.0980735e-32 * -446.85272 = 4.0654988e-29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010110010111100010111011001;
		b = 32'b01010110010000110111001101100010;
		correct = 32'b00111001100110111001001110001100;
		#400 //5.523274e-18 * 53725083000000.0 = 0.00029673835
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111010111010101101111111110;
		b = 32'b10110100111101010110111100011100;
		correct = 32'b10010100110101000011100100011101;
		#400 //4.6874664e-20 * -4.571565e-07 = -2.1429057e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010011011010011000000111001;
		b = 32'b11100100000001110000011011110010;
		correct = 32'b11101110111110100011010110111011;
		#400 //3886094.2 * -9.963244e+21 = -3.8718104e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100100011110001011110110000;
		b = 32'b11110100111011001001110110010010;
		correct = 32'b11110010000001000100000111101001;
		#400 //0.01746735 * -1.499729e+32 = -2.619629e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101111001100110111111100100;
		b = 32'b00110001010010110000100011111000;
		correct = 32'b00001111101101101100001011001101;
		#400 //6.0996185e-21 * 2.9545486e-09 = 1.802162e-29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110010001100001001001100101;
		b = 32'b10100111110100000001111110111000;
		correct = 32'b10111110101000010000011101111101;
		#400 //54445577000000.0 * -5.7765987e-15 = -0.31451026
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100100100010101100001100110;
		b = 32'b01011110110001111100000110010110;
		correct = 32'b00110011111000101101001101000000;
		#400 //1.4676125e-26 * 7.1969754e+18 = 1.0562371e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000000100011000010101010100;
		b = 32'b00110100010110100011100011111001;
		correct = 32'b01011100111110000001011111011000;
		#400 //2.7488104e+24 * 2.0323559e-07 = 5.586561e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111100111101001000111101011;
		b = 32'b11110010010011100001001101100100;
		correct = 32'b11111010011111110100101011011100;
		#400 //81187.836 * -4.0817506e+30 = -3.313885e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001101100111101110101001001;
		b = 32'b01000100110001100010110001000010;
		correct = 32'b00010111000010110011110000111111;
		#400 //2.8377598e-28 * 1585.383 = 4.4989364e-25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000100110101010000000110001;
		b = 32'b11001000110110001011011111110011;
		correct = 32'b01101010000000101110011001000101;
		#400 //-8.9135675e+19 * -443839.6 = 3.9561943e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101100001000010010101010010000;
		b = 32'b01001110100110110000000010110100;
		correct = 32'b00111011010000110010101001101101;
		#400 //2.2903103e-12 * 1300257300.0 = 0.0029779926
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110001010011001010100110111;
		b = 32'b00001000010001100100001110100000;
		correct = 32'b00101111000000110101011000110101;
		#400 //2.0020812e+23 * 5.966295e-34 = 1.1945007e-10
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100000101111011111010001011;
		b = 32'b11000111001011011011001111001010;
		correct = 32'b10011011110011011110110010101100;
		#400 //7.66113e-27 * -44467.79 = -3.406735e-22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111101011111101111101010110;
		b = 32'b10111010111111110001101010010011;
		correct = 32'b01100011001011110100000110111000;
		#400 //-1.6610679e+24 * -0.0019462876 = 3.2329157e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110000101110100100110111111;
		b = 32'b01001001011000110011110010110011;
		correct = 32'b01101000000001100100101001000011;
		#400 //2.7253636e+18 * 930763.2 = 2.536668e+24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110110100110000110001011001;
		b = 32'b01010101000101100000101111110000;
		correct = 32'b01011100011101110110011000100111;
		#400 //27014.174 * 10311126000000.0 = 2.7854655e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101010010110100011110000110;
		b = 32'b10000100010000010111000011011110;
		correct = 32'b00001010000110011001101010001100;
		#400 //-3252.4702 * -2.2738867e-36 = 7.395749e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110111001110110110101100110011;
		b = 32'b10010000010000011000001110010110;
		correct = 32'b11001000000011011010110000100111;
		#400 //3.8013038e+33 * -3.816391e-29 = -145072.61
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100011000011011011111011011;
		b = 32'b00101101011111110111001101010100;
		correct = 32'b10111010011000010011101111010011;
		#400 //-59170668.0 * 1.452068e-11 = -0.00085919834
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111100110001111101011001011;
		b = 32'b10101010111000100110111101111010;
		correct = 32'b10001011000001110101000000000101;
		#400 //6.4789406e-20 * -4.0223017e-13 = -2.6060254e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111110001010101100010100010;
		b = 32'b11101111100110100111110010110110;
		correct = 32'b11000111111011100010111011101001;
		#400 //1.2753201e-24 * -9.562292e+28 = -121949.82
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011111010000100010110111111;
		b = 32'b00100110101011100000010100011101;
		correct = 32'b01001011000111011110010000001011;
		#400 //8.569341e+21 * 1.2075061e-15 = 10347531.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110110101011101110101010011;
		b = 32'b11000100100001001100001100101010;
		correct = 32'b01100011110111011101001001010011;
		#400 //-7.7052824e+18 * -1062.0989 = 8.183772e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001001000101000101011111111;
		b = 32'b10100110111000110101001110011100;
		correct = 32'b11011000100100000101011001010110;
		#400 //8.048737e+29 * -1.5773952e-15 = -1269603900000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000010110111101000011110111;
		b = 32'b11101110010001111111011110010110;
		correct = 32'b01000111001010111011010000000111;
		#400 //-2.8410587e-24 * -1.5471707e+28 = 43956.027
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111111100011100001000111110;
		b = 32'b01000011111100101100101001010110;
		correct = 32'b11101100011001010100100010110011;
		#400 //-2.2833469e+24 * 485.58075 = -1.1087493e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110111000010011111001100110;
		b = 32'b10000001000010100001101000110100;
		correct = 32'b10011000011100110000010101100010;
		#400 //123829060000000.0 * -2.5365397e-38 = -3.1409732e-24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101101000010100011011111010;
		b = 32'b01001111111111010111010001001010;
		correct = 32'b11000110000111111010110001101000;
		#400 //-1.2016092e-06 * 8504513500.0 = -10219.102
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111000101111010101111000100;
		b = 32'b11001101100000111000010000010110;
		correct = 32'b01111101000110111101011001001110;
		#400 //-4.693989e+28 * -275808960.0 = 1.2946442e+37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011110010000001010100110001;
		b = 32'b10110011001111100011101110100000;
		correct = 32'b10100111100101001010111001010100;
		#400 //9.3170804e-08 * -4.429205e-08 = -4.126726e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110000011010101011001111111;
		b = 32'b10111110000100101100111100101010;
		correct = 32'b00101100101000100001101101101001;
		#400 //-3.2136512e-11 * -0.1433684 = 4.60736e-12
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010101001000010010111010010;
		b = 32'b00000100100011010101100100101001;
		correct = 32'b10000111101101010100010000000000;
		#400 //-82.07387 * 3.323082e-36 = -2.727382e-34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100110100101110001110111100;
		b = 32'b00000000010101010100110011000110;
		correct = 32'b00001101100011001000100110111000;
		#400 //110566880.0 * 7.833558e-39 = 8.661321e-31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001001111001100101100010110;
		b = 32'b00111000010000100000100110010001;
		correct = 32'b10010010000011110001100011110101;
		#400 //-9.760385e-24 * 4.6262114e-05 = -4.5153606e-28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111000111101010011011100000;
		b = 32'b11100011011001101111010101100001;
		correct = 32'b01011011000011110010000111111111;
		#400 //-9.4563875e-06 * -4.2604326e+21 = 4.02883e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110011011010110100100101110;
		b = 32'b10100000000111001010010101010101;
		correct = 32'b11000111000100010100010101101100;
		#400 //2.8028527e+23 * -1.3268418e-19 = -37189.42
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010010100111100110000010001;
		b = 32'b00011001101100000010010110011111;
		correct = 32'b10000100100100011011101101101100;
		#400 //-1.8811364e-13 * 1.8213169e-23 = -3.4261456e-36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100010101010100110101011110;
		b = 32'b10000010011010001110110000000011;
		correct = 32'b10000111010000100001001011000011;
		#400 //853.20886 * -1.71124e-37 = -1.4600451e-34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101001101111100110001000100;
		b = 32'b10011111100101001010101110000001;
		correct = 32'b10000101010101010111101001110011;
		#400 //1.5941928e-16 * -6.296417e-20 = -1.0037702e-35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110111111100111010011010001;
		b = 32'b00010011111101101101011111000101;
		correct = 32'b11010011011101010101101010111001;
		#400 //-1.6911523e+38 * 6.2311896e-27 = -1053789060000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011101101001000111000011010;
		b = 32'b00110001010011010010101000100111;
		correct = 32'b01100101100100001011001110000110;
		#400 //2.8610095e+31 * 2.9855387e-09 = 8.541655e+22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110000000010100111100101111;
		b = 32'b10010111001111111010011111011010;
		correct = 32'b10111101110000011001110110111010;
		#400 //1.5266149e+23 * -6.1927287e-25 = -0.09453912
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101001101000001000010101111;
		b = 32'b01010111011111110010110111110100;
		correct = 32'b10111101001100110111110011110001;
		#400 //-1.5618164e-16 * 280572830000000.0 = -0.043820325
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101001000000100011110100000;
		b = 32'b00111011110100010000010010001001;
		correct = 32'b00111001100000101101110101010001;
		#400 //0.039130807 * 0.0063787145 = 0.00024960426
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110101001001111010001011111;
		b = 32'b11010101101110000001101111101101;
		correct = 32'b10110100111011010100001101000110;
		#400 //1.7465245e-20 * -25303760000000.0 = -4.4193638e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101111001010001100010001011;
		b = 32'b10010110100100010110111101111000;
		correct = 32'b00101101000000100010011010101000;
		#400 //-31486697000000.0 * -2.349636e-25 = 7.398228e-12
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010111010011001111000110101;
		b = 32'b00011001100000010000100000111110;
		correct = 32'b01000100111010111000000001111100;
		#400 //1.4121341e+26 * 1.3341616e-23 = 1884.0151
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101110001100000101010000000;
		b = 32'b00101111011001100011010101101110;
		correct = 32'b11100101101100100001011011000100;
		#400 //-5.0209362e+32 * 2.093736e-10 = -1.0512515e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001101101011110010100011110;
		b = 32'b10011011001011011111010100101000;
		correct = 32'b00000101011101110011010000001100;
		#400 //-8.07776e-14 * -1.4389439e-22 = 1.1623444e-35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001000110100010110100111111;
		b = 32'b10000000010010011100001010100000;
		correct = 32'b00101001101100011011000001110110;
		#400 //-1.1649265e+25 * -6.77381e-39 = 7.89099e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011110011001110000110001110;
		b = 32'b10100001000000010010110101110011;
		correct = 32'b11001101010011101100010000010000;
		#400 //4.9537204e+26 * -4.376705e-19 = -216809730.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011011000011110101000101000;
		b = 32'b11010111110011001110011000110001;
		correct = 32'b01011011101101001101000110111011;
		#400 //-225.91467 * -450578070000000.0 = 1.0179219e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111011100010101010011001011;
		b = 32'b01010110000100000001110111001011;
		correct = 32'b01100110000001111101101111001000;
		#400 //4048866000.0 * 39614410000000.0 = 1.6039343e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110010101110011001100110111;
		b = 32'b10111000111011111101100011101000;
		correct = 32'b10111111110010011001111100100111;
		#400 //13772.804 * -0.0001143681 = -1.5751694
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110111110011100111011001111;
		b = 32'b10011110010010101001110111101100;
		correct = 32'b10100101110001011011011101001001;
		#400 //31975.404 * -1.07264484e-20 = -3.4298251e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011100011011010011111010111;
		b = 32'b01010110101001001100000000001101;
		correct = 32'b11110010101101100101001110010110;
		#400 //-7.974503e+16 * 90572380000000.0 = -7.222697e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011011010010000110000111111;
		b = 32'b11011001100000111010110001001110;
		correct = 32'b00110101011011111011110000111111;
		#400 //-1.9277265e-22 * -4632834000000000.0 = 8.930837e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100011010100000010101100010;
		b = 32'b00011101011110011101110110110100;
		correct = 32'b00011010011001000110100111101000;
		#400 //0.01428351 * 3.3069493e-21 = 4.7234845e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011011011101011011110100010;
		b = 32'b00010000010001011001101110011000;
		correct = 32'b10000100001110000100010001100111;
		#400 //-5.5580706e-08 * 3.8971265e-29 = -2.1660505e-36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110010001101001100001100100;
		b = 32'b00110110010110100011101110001111;
		correct = 32'b00010101001010010100101111111001;
		#400 //1.0513546e-20 * 3.25192e-06 = 3.418921e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001001011101110001011010011;
		b = 32'b10111011001011110011001010110001;
		correct = 32'b01100100111011110101111101011111;
		#400 //-1.3214015e+25 * -0.0026733095 = 3.5325152e+22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001101101000111101011110101;
		b = 32'b10011001100000001010010100011001;
		correct = 32'b01001011101101010110001110111111;
		#400 //-1.7873903e+30 * -1.3301572e-23 = 23775102.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000011101010101011001000010;
		b = 32'b11110111011011100111010011100010;
		correct = 32'b01010000011001001000011000110101;
		#400 //-3.1709057e-24 * -4.836474e+33 = 15336003000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101000100011001000110100110;
		b = 32'b00100000100010011011101000110011;
		correct = 32'b10011110000111001010000110100101;
		#400 //-0.03553929 * 2.333192e-19 = -8.2919985e-21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001010000000001011100011101;
		b = 32'b01100111010000110000001100100100;
		correct = 32'b11010001000100100101001111110110;
		#400 //-4.2652612e-14 * 9.209194e+23 = -39279616000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110001011111101101100001001;
		b = 32'b00111010010101110110010001100000;
		correct = 32'b00110001000100111111010111101000;
		#400 //2.6204527e-06 * 0.0008216556 = 2.1531097e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011010010110010100110010000;
		b = 32'b01011111111011000011100110110011;
		correct = 32'b01001011101110110111100000011011;
		#400 //7.2177767e-13 * 3.4043666e+19 = 24571958.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001110011111011101110000000;
		b = 32'b11000010101110110111010000011110;
		correct = 32'b10111101000110000001110000110000;
		#400 //0.00039621815 * -93.72679 = -0.037136257
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101100001100100011100110110010;
		b = 32'b00100000111000111001001000010001;
		correct = 32'b00001101100111100110111011011010;
		#400 //2.5327349e-12 * 3.8551954e-19 = 9.764188e-31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000110110000001100011011011;
		b = 32'b11011110000010111010101001001001;
		correct = 32'b01100111011010111100101001111010;
		#400 //-442566.84 * -2.5159841e+18 = 1.11349116e+24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101010000010000111111111001;
		b = 32'b11011110101111001011100110101100;
		correct = 32'b01001100100011100101001111000001;
		#400 //-1.09743265e-11 * -6.799545e+18 = 74620424.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111010111110111101110000101;
		b = 32'b11010111100010010100010001000110;
		correct = 32'b11011111011011111010100101101000;
		#400 //57211.52 * -301852650000000.0 = -1.7269449e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011001111010000100010111100;
		b = 32'b11110010110000100100010000110100;
		correct = 32'b01011110100011110111001011111011;
		#400 //-6.715841e-13 * -7.6956857e+30 = 5.1683e+18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011000100011001010010010010;
		b = 32'b00111111011011111001001010000010;
		correct = 32'b01010011000010000011110100000101;
		#400 //625262850000.0 * 0.9358293 = 585139300000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101100110011100111000000110;
		b = 32'b10011001101100110111010001100010;
		correct = 32'b01001111110101111010000111110101;
		#400 //-3.8994144e+32 * -1.8555173e-23 = 7235431000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101010100100110001000101110;
		b = 32'b11110111001111110111010010001011;
		correct = 32'b11001101000111010101011100000111;
		#400 //4.2486612e-26 * -3.8831737e+33 = -164982900.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100010001010010101010000010;
		b = 32'b00100101001100010001011111001111;
		correct = 32'b00100010000010000110010010111010;
		#400 //0.01203406 * 1.536037e-16 = 1.8484761e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110010110001111010101101011;
		b = 32'b00000110011101011111000100110000;
		correct = 32'b10111101010100000110111101000111;
		#400 //-1.1001111e+33 * 4.6256575e-35 = -0.050887372
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000011101110001100001001100;
		b = 32'b00000000111111010010010101100000;
		correct = 32'b00010001111101000101011100010110;
		#400 //16582259000.0 * 2.3247788e-38 = 3.8550083e-28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000000010011010111101101100;
		b = 32'b01010110110001010010000111101011;
		correct = 32'b01101111010101000000110001111000;
		#400 //605546100000000.0 * 108374730000000.0 = 6.5625896e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000011011000110011111111100;
		b = 32'b00100101111100111011010011010011;
		correct = 32'b10111110111000010000110110110000;
		#400 //-1039725400000000.0 * 4.2276312e-16 = -0.43955755
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110010110110010111100100100;
		b = 32'b00101100110001000011001011001111;
		correct = 32'b11010011101001111111101110011000;
		#400 //-2.5876696e+23 * 5.576296e-12 = -1442961200000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001100010001110001111000100;
		b = 32'b00111100001101111000010110101010;
		correct = 32'b11100110010001000100010010010101;
		#400 //-2.0686188e+25 * 0.011201302 = -2.3171224e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110010111001101100000000100;
		b = 32'b01000111001101101100100011101010;
		correct = 32'b10111110000111011010111011100101;
		#400 //-3.2908292e-06 * 46792.914 = -0.15398748
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111100111110110011011110010;
		b = 32'b11011111011011111100011011011001;
		correct = 32'b11000111100101010100110011101101;
		#400 //4.424298e-15 * -1.7277736e+19 = -76441.85
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111110111000001011011101001;
		b = 32'b10110010111001100011000110101000;
		correct = 32'b01100011010001011110011101000110;
		#400 //-1.362288e+29 * -2.6798105e-08 = 3.6506736e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001100101011001011100100011;
		b = 32'b10110111100000011001000001111010;
		correct = 32'b11101001100101110110101100101010;
		#400 //1.4814713e+30 * -1.5445275e-05 = -2.2881733e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010000101001111110001001001;
		b = 32'b10000110100000001000010011001011;
		correct = 32'b00000001000101011001011011011001;
		#400 //-0.00056833454 * -4.834337e-35 = 2.7475206e-38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111000001101110001010110000;
		b = 32'b01010100101111111011101001001101;
		correct = 32'b11110100010010100000101010010101;
		#400 //-9.719524e+18 * 6587715000000.0 = -6.4029455e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100111110110001111000101000;
		b = 32'b00110010110100101101011010110000;
		correct = 32'b00111000010011101101000101010101;
		#400 //2008.9424 * 2.4544846e-08 = 4.9309183e-05
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110111000101011001111011000;
		b = 32'b01100010001010101010110100010000;
		correct = 32'b01011001100101110010010010101111;
		#400 //6.7562614e-06 * 7.8710424e+20 = 5317882000000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011001011010110011011110101;
		b = 32'b10110100010000001100011000010111;
		correct = 32'b11010000000000101001001101100101;
		#400 //4.8808373e+16 * -1.7953458e-07 = -8762791000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100000110000110100111111101;
		b = 32'b01001100100001100001101101001000;
		correct = 32'b10111001000111111010111101110001;
		#400 //-2.1659334e-12 * 70310460.0 = -0.00015228779
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100000011101000001101110001;
		b = 32'b11100010010011100000100011011111;
		correct = 32'b11101110111001010110010101101010;
		#400 //37359044.0 * -9.501671e+20 = -3.5497335e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011111110110100010100100011;
		b = 32'b01111000011001001001001010101000;
		correct = 32'b01001100111000000101100110000101;
		#400 //6.3429482e-27 * 1.8544035e+34 = 117623850.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101111011100111000010100000;
		b = 32'b01010011001100111100100100110000;
		correct = 32'b11011001101001110111010000100011;
		#400 //-7630.078 * 772174500000.0 = -5891752000000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110000011110110101011010101;
		b = 32'b01000011001000100011101000001100;
		correct = 32'b10101001101101011100010000111111;
		#400 //-4.9757876e-16 * 162.22675 = -8.072058e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100001010000011100100000010;
		b = 32'b00001001010011010111100101101100;
		correct = 32'b10100110000001110000010101110001;
		#400 //-1.894019e+17 * 2.473307e-33 = -4.684491e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111100010110100001100000100;
		b = 32'b00110101010100010101110010110000;
		correct = 32'b10001101011000111100100001000100;
		#400 //-8.999582e-25 * 7.7993445e-07 = -7.0190837e-31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001010001110111111111001111;
		b = 32'b11011100011110001100000010001000;
		correct = 32'b00011110010000011101100111011010;
		#400 //-3.6642226e-38 * -2.8006994e+17 = 1.02623856e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011001001001011001111111010;
		b = 32'b11010000110100001001010001100101;
		correct = 32'b00100100100001100011000110110100;
		#400 //-2.0788445e-27 * -27995089000.0 = 5.819744e-17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100011111100010111100100001;
		b = 32'b00110010011101101110010010001101;
		correct = 32'b11010111011101010010010000111000;
		#400 //-1.8755476e+22 * 1.4371051e-08 = -269535900000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010101100101010001000001100;
		b = 32'b10001010011101001110010101101101;
		correct = 32'b00100101101010101110001010001010;
		#400 //-2.514036e+16 * -1.1791323e-32 = 2.9643808e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011110110011110101010011101;
		b = 32'b10110100111001001101111011111000;
		correct = 32'b00100001010000101101001011000000;
		#400 //-1.5483896e-12 * -4.263054e-07 = 6.600868e-19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100100110011101110101100010;
		b = 32'b00001111001010100101011011111011;
		correct = 32'b00101100010011001100001010010101;
		#400 //3.4647268e+17 * 8.398399e-30 = 2.9098158e-12
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011001010110001110001011111;
		b = 32'b11000011101111101101110011001101;
		correct = 32'b11010111011111110010010101001000;
		#400 //734915400000.0 * -381.725 = -280535590000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001101001111100010010101101;
		b = 32'b01001000001011110010100101010000;
		correct = 32'b11011010011001011001010100001010;
		#400 //-90069900000.0 * 179365.25 = -1.615541e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111100100011111001100101000010;
		b = 32'b00000010110100111110110001001010;
		correct = 32'b00111111111011011011111110111000;
		#400 //5.964855e+36 * 3.1139287e-37 = 1.8574133
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110000111111110110010101010;
		b = 32'b00111111011000011000010011011000;
		correct = 32'b10101110000011001110000111111110;
		#400 //-3.6362614e-11 * 0.8809333 = -3.2033036e-11
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101001011101111000010011110;
		b = 32'b10011101001101110010001001010000;
		correct = 32'b11010010111110100100101011100111;
		#400 //2.2176268e+32 * -2.4237587e-21 = -537499240000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010111101111111110011000100;
		b = 32'b01100011001001000101010100111110;
		correct = 32'b01100110100111110011000010000001;
		#400 //123.99368 * 3.0314084e+21 = 3.758755e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011011010100000111011110011;
		b = 32'b00001100000100010110010110111101;
		correct = 32'b00110000000001001110111101111100;
		#400 //4.3176153e+21 * 1.120101e-31 = 4.836165e-10
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110011101001110000110000110;
		b = 32'b01100111100010000101000001011111;
		correct = 32'b10110110100000100110010010110001;
		#400 //-3.0183908e-30 * 1.2874489e+24 = -3.886024e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111000110011110100001111111;
		b = 32'b00000111001111110010010000111010;
		correct = 32'b00001110111001011101010001111101;
		#400 //39400.496 * 1.4379889e-34 = 5.6657477e-30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001000000101000001011001000;
		b = 32'b11111111000110101100001110111000;
		correct = 32'b01001000100111011100110011100111;
		#400 //-1.5709674e-33 * -2.0571734e+38 = 323175.22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011010001101110110000101010;
		b = 32'b11010000111000110111010110001101;
		correct = 32'b11110100101100001011111011000001;
		#400 //3.6694727e+21 * -30529055000.0 = -1.1202554e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001100010001010001100001110;
		b = 32'b10001000100100000111000100100011;
		correct = 32'b11000010100110100011000000110101;
		#400 //8.868244e+34 * -8.693283e-34 = -77.094154
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110101110100011100100100101;
		b = 32'b00011001101100010100001111001111;
		correct = 32'b00110001000000001111001011010110;
		#400 //102377300000000.0 * 1.8328759e-23 = 1.8764488e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111010100101110011001110111;
		b = 32'b00111100010001110001010000100101;
		correct = 32'b00010100001001000000000110111111;
		#400 //6.8145547e-25 * 0.012150799 = 8.2802284e-27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100001110011000110100000011;
		b = 32'b00110100110011011100001010110101;
		correct = 32'b10000001100101010010001100001011;
		#400 //-1.4294316e-31 * 3.8325894e-07 = -5.478424e-38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000010110011000000000101110111;
		b = 32'b11111100000011010011011011001001;
		correct = 32'b00111111011000010001000011101110;
		#400 //-2.9975947e-37 * -2.9329e+36 = 0.8791646
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100000100111010001001000111;
		b = 32'b01001000111010011001101111101111;
		correct = 32'b01110101100001101011100010100000;
		#400 //7.139137e+26 * 478431.47 = 3.415588e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111000001111110000101101000100;
		b = 32'b10110001100010010111111011011110;
		correct = 32'b10101010010011010011011101101001;
		#400 //4.554844e-05 * -4.001648e-09 = -1.8226882e-13
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000110001110110010011000001;
		b = 32'b01101100110100001011110100001110;
		correct = 32'b01101110001000101001010100011101;
		#400 //6.231049 * 2.0187948e+27 = 1.257921e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100011101000001001111110110;
		b = 32'b10111011101011111000110101110100;
		correct = 32'b00111000101001110110000010000011;
		#400 //-0.014897337 * -0.0053574387 = 7.981157e-05
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011101000010000010001001011;
		b = 32'b10001000101100001001110000010000;
		correct = 32'b10001100110111100010101000111000;
		#400 //322.03354 * -1.0629305e-33 = -3.4229925e-31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100101110111000000111000001;
		b = 32'b00100011111100100010100000100001;
		correct = 32'b00110001001100010101111000001101;
		#400 //98307590.0 * 2.6254688e-17 = 2.5810352e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001010001000111101001011110;
		b = 32'b10100001100000011100000111111000;
		correct = 32'b10010011010001110010110100010000;
		#400 //2.8591312e-09 * -8.792723e-19 = -2.5139549e-27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000001101011000011010100100;
		b = 32'b00101000010101101000111000110001;
		correct = 32'b11011001000110000010001101100001;
		#400 //-2.2471823e+29 * 1.1910219e-14 = -2676443500000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100110011010101010100000010;
		b = 32'b00011010111100001110001011110110;
		correct = 32'b11000000010000010011010110111100;
		#400 //-3.0301664e+22 * 9.962835e-23 = -3.0189047
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010110001101000010001011001;
		b = 32'b01111111011101111011001010001000;
		correct = 32'b11101010110000000001010000100011;
		#400 //-3.52637e-13 * 3.292463e+38 = -1.16104425e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101000101001110100010101000;
		b = 32'b10000011010101101000110010011010;
		correct = 32'b00100000111110011001100010001010;
		#400 //-6.706257e+17 * -6.305035e-37 = 4.2283183e-19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101101111111111011100010101;
		b = 32'b10101110010000110110101110110011;
		correct = 32'b11001100100100101000100111110111;
		#400 //1.7290685e+18 * -4.4433523e-11 = -76828600.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111011100011010111111100000;
		b = 32'b10010000000100110011000101101101;
		correct = 32'b00100000000010101111011010100111;
		#400 //-4054835200.0 * -2.9028715e-29 = 1.1770665e-19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010111100101010101110001110;
		b = 32'b01010101001100010101100000101000;
		correct = 32'b00110000101010000001110000101110;
		#400 //1.00366016e-22 * 12187012000000.0 = 1.2231618e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111110110110010000001111001;
		b = 32'b01110111101000100000010000101011;
		correct = 32'b01111111110110110010000001111001;
		#400 //nan * 6.572161e+33 = nan
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111110111010110110010100100;
		b = 32'b01101101001000110010101011011000;
		correct = 32'b00111101100011010010000100111011;
		#400 //2.183413e-29 * 3.1561157e+27 = 0.06891104
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010011110110001000011001001;
		b = 32'b01100111110010111101010111000101;
		correct = 32'b11100010110001111110011111110110;
		#400 //-0.00095773913 * 1.9251675e+24 = -1.8438083e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101011110000010111011101001;
		b = 32'b10000101010010100010110100001001;
		correct = 32'b00011011010001000000000010101101;
		#400 //-17055023000000.0 * -9.506266e-36 = 1.6212958e-22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000110001101000100011011000;
		b = 32'b11111011001101011111101110111110;
		correct = 32'b10111100100011010010000111111100;
		#400 //1.8232519e-38 * -9.449117e+35 = -0.01722812
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110001101100110100010101011;
		b = 32'b11100111111000001111101110010110;
		correct = 32'b10110110101000000100111011011001;
		#400 //2.2483628e-30 * -2.124902e+24 = -4.7775507e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000100101011111100110010001;
		b = 32'b00011111100010010110101000111101;
		correct = 32'b10000000101000010000000110010111;
		#400 //-2.540673e-19 * 5.8197513e-20 = -1.4786085e-38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001011110001010011110010110;
		b = 32'b10100001001110010011111100001001;
		correct = 32'b01010011001100111110111001010101;
		#400 //-1.2312781e+30 * -6.2763864e-19 = 772797700000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000001100111011010011111000;
		b = 32'b10110111010110011000011101001101;
		correct = 32'b01000000000110001011001101100001;
		#400 //-184019.88 * -1.296571e-05 = 2.3859484
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000010001000111001000001101101;
		b = 32'b01001010100001111101101101111111;
		correct = 32'b10001101001011011001101011001110;
		#400 //-1.2016797e-37 * 4451775.5 = -5.349608e-31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111011111100110111100000011;
		b = 32'b10000111111101001010010001000110;
		correct = 32'b10010111111100110010010100010100;
		#400 //4268688100.0 * -3.680959e-34 = -1.5712867e-24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010011100110011001111011010;
		b = 32'b01101010011100110011011110011100;
		correct = 32'b01101101011001110000111100001100;
		#400 //60.800636 * 7.3507896e+25 = 4.4693267e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111110001100010111000001110;
		b = 32'b11011101100011110100001000111010;
		correct = 32'b01101101110111011100110111111101;
		#400 //-6649814000.0 * -1.2903596e+18 = 8.5806515e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011011101101111000111100001;
		b = 32'b01001011110110110001101100100100;
		correct = 32'b00011111110100110101101100011010;
		#400 //3.116882e-27 * 28718664.0 = 8.951269e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011111100011110111110101101;
		b = 32'b10111110101000111100101010111101;
		correct = 32'b10001011000110101100101100110101;
		#400 //9.319045e-32 * -0.31990615 = -2.9812197e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001011101100001111000011110;
		b = 32'b01001010101011100110000001000101;
		correct = 32'b11101100101001111010010100000110;
		#400 //-2.8375433e+20 * 5713954.5 = -1.6213593e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110101011000011001101100000;
		b = 32'b00000101111101010110000000011111;
		correct = 32'b00010101001001010000110111010011;
		#400 //1444524000.0 * 2.3074999e-35 = 3.333239e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101000111101010001111111110;
		b = 32'b00100000010011001111000011111101;
		correct = 32'b10011101111111100000000000001010;
		#400 //-0.038730614 * 1.7359208e-19 = -6.723328e-21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111000001110010010111001111;
		b = 32'b00010011010001010010010101101110;
		correct = 32'b00001010110100000010011110110110;
		#400 //8.05543e-06 * 2.488335e-27 = 2.0044609e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100101110001100111100111000;
		b = 32'b01101101100110100101000110000010;
		correct = 32'b01110010110111101100111011111110;
		#400 //1478.4756 * 5.9699036e+27 = 8.8263565e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101010011111011110010000100;
		b = 32'b00010101111011101110111111011000;
		correct = 32'b00111011110000011110001111100011;
		#400 //6.131296e+22 * 9.650584e-26 = 0.005917059
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100100100001001101010001011;
		b = 32'b00001010011110010001001100100111;
		correct = 32'b10010111100011001011000100100011;
		#400 //-75813976.0 * 1.1992516e-32 = -9.092004e-25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101000111101100101001110011;
		b = 32'b00100010011011110010110010101010;
		correct = 32'b10010000000101000101101010110110;
		#400 //-9.026213e-12 * 3.2414185e-18 = -2.9257735e-29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010011111111101010100100101;
		b = 32'b10111100010001100011111100001001;
		correct = 32'b00101111010001100001110111011001;
		#400 //-1.4891417e-08 * -0.01209999 = 1.8018599e-10
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000010001100101000010000111;
		b = 32'b10111010011000010110010000110100;
		correct = 32'b00001011001011101001101001100110;
		#400 //-3.911065e-29 * -0.0008598 = 3.3627338e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010001011010010101110110100;
		b = 32'b01100010001111001011000100100010;
		correct = 32'b10101100111111110100011111010101;
		#400 //-8.337867e-33 * 8.701879e+20 = -7.255511e-12
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010000010000111010011111000;
		b = 32'b11011100110010001001011100101011;
		correct = 32'b01001111010101011101011111101011;
		#400 //-7.9428375e-09 * -4.5168965e+17 = 3587697400.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110010001001100111011111001;
		b = 32'b11001110100001000110001001011010;
		correct = 32'b11100101010010111000110010101010;
		#400 //54098305000000.0 * -1110519000.0 = -6.00772e+22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100001000110010010100010110;
		b = 32'b01010110110101011011001010000101;
		correct = 32'b01111011100010000010111110100000;
		#400 //1.2037966e+22 * 117481360000000.0 = 1.4142366e+36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111011001100101011110001100;
		b = 32'b11001001011011111101110110000110;
		correct = 32'b11111001010101111101001100001110;
		#400 //7.128739e+28 * -982488.4 = -7.0039033e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111110011010111001011110000;
		b = 32'b10101000111001000111010110000000;
		correct = 32'b10101001001101110101100010101010;
		#400 //1.6050701 * -2.5364042e-14 = -4.0711067e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111100110000101110010111100;
		b = 32'b00101111010100100011111110011000;
		correct = 32'b00000111011110100100001111010111;
		#400 //9.846179e-25 * 1.9121982e-10 = 1.8827846e-34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101011110101010101001000101;
		b = 32'b01110101011101110001000000110100;
		correct = 32'b11011011011100011110101000100110;
		#400 //-2.1741733e-16 * 3.1318993e+32 = -6.809292e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111010100011111011110110011100;
		b = 32'b00110110111011001111111100001001;
		correct = 32'b11110010000001010001000111111111;
		#400 //-3.731721e+35 * 7.063038e-06 = -2.6357288e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110111111000000010000010000;
		b = 32'b00010001000100111101000100111010;
		correct = 32'b00001000100100011000010001001110;
		#400 //7.510658e-06 * 1.1660728e-28 = 8.757975e-34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101001100000001000010001010;
		b = 32'b10111000111110100001110111000001;
		correct = 32'b01110110101011000000010010011101;
		#400 //-1.4626875e+37 * -0.00011926471 = 1.74447e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110101110011010101100111000;
		b = 32'b10111010000000110010110000001000;
		correct = 32'b11111001001111100100010100011010;
		#400 //1.233981e+38 * -0.00050038146 = -6.174612e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101000111111111010100110001;
		b = 32'b01001001000101000001100110010011;
		correct = 32'b10100110101110010001001101110110;
		#400 //-2.1170236e-21 * 606617.2 = -1.2842229e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101110110011101101011100010;
		b = 32'b01111000001000010001000100011110;
		correct = 32'b11110110100010010001000100111001;
		#400 //-0.10637452 * 1.3067296e+34 = -1.3900273e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101110100110001011001000100;
		b = 32'b11001111110101001001100101011010;
		correct = 32'b01111110001011110100110011100011;
		#400 //-8.166032e+27 * -7133639700.0 = 5.825353e+37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010010100010110000101100101;
		b = 32'b00100111110100110000100110000100;
		correct = 32'b00011010101011001001101100001111;
		#400 //1.2187546e-08 * 5.857458e-15 = 7.1388043e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111011001110010010111101101;
		b = 32'b01001000010110011101010100101110;
		correct = 32'b01101000010001001010111110100010;
		#400 //1.6655979e+19 * 223060.72 = 3.7152947e+24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110111110011100100100000010;
		b = 32'b00011010110101010010110110100101;
		correct = 32'b11010010010100000000000011001000;
		#400 //-2.5331227e+33 * 8.816848e-23 = -223341580000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010001111101001000001101110;
		b = 32'b01011111010011010001100101110101;
		correct = 32'b11100010000110001010110010011011;
		#400 //-47.641045 * 1.4778972e+19 = -7.0408566e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111111101101001001010100111;
		b = 32'b10110000101001100011001110011101;
		correct = 32'b00011001001000000001010011001111;
		#400 //-6.8437717e-15 * -1.2092759e-09 = 8.276008e-24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000110110110010101010100111;
		b = 32'b01110000001101111010111010111001;
		correct = 32'b01010001100111010100000100010011;
		#400 //3.7128268e-19 * 2.2738793e+29 = 84425200000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110001010010000101110110011;
		b = 32'b11101011011100010011011100101111;
		correct = 32'b01101010000111110100100001110100;
		#400 //-0.16508369 * -2.9161172e+26 = 4.814034e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100111110100110111100010010;
		b = 32'b01001010011001101100111111111111;
		correct = 32'b10111111111000011100101101000011;
		#400 //-4.6646943e-07 * 3781631.8 = -1.7640156
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010000111011010101010011000;
		b = 32'b11001100011001011100111011000001;
		correct = 32'b00011111000011011000100011110000;
		#400 //-4.975074e-28 * -60242692.0 = 2.9971183e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100101000001010110101101001;
		b = 32'b01111000000011011011000001100111;
		correct = 32'b01101101001100011101110001110101;
		#400 //2.9928495e-07 * 1.1495183e+34 = 3.4403352e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111010101001101010101100011001;
		b = 32'b00010001011001111100001100100000;
		correct = 32'b11001100100101101110001101101101;
		#400 //-4.3269578e+35 * 1.8282814e-28 = -79108970.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100001011110100001100010100;
		b = 32'b10111001101000111110101101110001;
		correct = 32'b00000110011000000111000111001011;
		#400 //-1.3501695e-31 * -0.000312652 = 4.221332e-35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111001010010011110100101001;
		b = 32'b11011000111001100001111001100001;
		correct = 32'b10111000100110000010000100001000;
		#400 //3.5837733e-20 * -2024145200000000.0 = -7.254077e-05
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000000111110000001111010111;
		b = 32'b00100000100000010111000111111001;
		correct = 32'b00101001001000001100111101110101;
		#400 //162831.36 * 2.192887e-19 = 3.5707077e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101001011110101011110001110;
		b = 32'b01001100000001110001101100000111;
		correct = 32'b00101001101110010001001101011110;
		#400 //2.3206322e-21 * 35417116.0 = 8.21901e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001000010011111000111001000;
		b = 32'b10101110100101111101101010011001;
		correct = 32'b01000000001000111010011011001111;
		#400 //-37029183000.0 * -6.905516e-11 = 2.5570562
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011001100011000011010100110;
		b = 32'b00001010001011011101111001011010;
		correct = 32'b10101101111100010010010001011111;
		#400 //-3.2747761e+21 * 8.371467e-33 = -2.741468e-11
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000100001001100110100011011;
		b = 32'b00101010001010110111101001100110;
		correct = 32'b01010011001100011110100011111111;
		#400 //5.017087e+24 * 1.5230316e-13 = 764118240000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110000100111010110101011010;
		b = 32'b10000110011111100100001000110011;
		correct = 32'b00110101000100101010110000101111;
		#400 //-1.1425966e+28 * -4.7820726e-35 = 5.46398e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101001011010110110001010101;
		b = 32'b11100000010011100111100011010001;
		correct = 32'b10110110000010111101111100000101;
		#400 //3.502253e-26 * -5.9511485e+19 = -2.0842429e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000110010000010000101100011;
		b = 32'b01010010011100011011101001100110;
		correct = 32'b00011011101111001111100100100110;
		#400 //1.2044911e-33 * 259553590000.0 = 3.1263e-22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000101100101011111000100010;
		b = 32'b11100000001001111010101101111110;
		correct = 32'b11100001011010100010001110001010;
		#400 //5.5857096 * -4.8327556e+19 = -2.6994369e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110100000010100111000110100;
		b = 32'b00000011110110011001110111110111;
		correct = 32'b10100010110110111101011000101000;
		#400 //-4.658721e+18 * 1.2790381e-36 = -5.9586816e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011110000010110011100100000;
		b = 32'b00101010010001011000111000111011;
		correct = 32'b00111110100101010011111111001111;
		#400 //1661317700000.0 * 1.7546461e-13 = 0.29150245
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011001001100101100111111010;
		b = 32'b10100100000000101001010000011000;
		correct = 32'b01011111101010011011001111011001;
		#400 //-8.637462e+35 * -2.8314697e-17 = 2.4456712e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101101001110111110111111000101;
		b = 32'b00100110110001101111110111011001;
		correct = 32'b00010100100100100001010111001110;
		#400 //1.0682959e-11 * 1.3807815e-15 = 1.4750833e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111000110011001001101101000101;
		b = 32'b00101000100000011010001000101111;
		correct = 32'b11100001110011110011011110111011;
		#400 //-3.3199306e+34 * 1.4392213e-14 = -4.7781148e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010101011010011110100001101;
		b = 32'b11001011010000111110011010110101;
		correct = 32'b10010110100001001001000110100000;
		#400 //1.6682259e-32 * -12838581.0 = -2.1417652e-25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001110100001111000011101111;
		b = 32'b01000101001010110010101011100011;
		correct = 32'b01110111100010111011001111110000;
		#400 //2.0692529e+30 * 2738.6804 = 5.667022e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010100101101011100001101001;
		b = 32'b11101110010100101001111110101101;
		correct = 32'b10111001011110000000001010010001;
		#400 //1.4513842e-32 * -1.6296222e+28 = -0.00023652079
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101101001010010100101110100011;
		b = 32'b10011101000110110000101010110011;
		correct = 32'b10001010110011010000111110111110;
		#400 //9.6233325e-12 * -2.051961e-21 = -1.9746703e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110100000001001111011001000;
		b = 32'b01001001000010100001010101000111;
		correct = 32'b01000000000010101100000010010001;
		#400 //3.833182e-06 * 565588.44 = 2.1680033
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001111000011000000000110111;
		b = 32'b00101110101110110100001111001010;
		correct = 32'b11000001001001001111010001011111;
		#400 //-121064840000.0 * 8.515817e-11 = -10.309661
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110011011011010111011001000;
		b = 32'b00011001100101110101111101100110;
		correct = 32'b11001000100011001000101010101011;
		#400 //-1.8389811e+28 * 1.5651565e-23 = -287829.34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010111100110001011011101001;
		b = 32'b00111100001110011000111101011010;
		correct = 32'b00100111101100000011001110101110;
		#400 //4.3181368e-13 * 0.011325682 = 4.8905844e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100101100010111001100010010;
		b = 32'b00110000001001111000110001001011;
		correct = 32'b11011101011010000100011010011111;
		#400 //-1.7161862e+27 * 6.0953614e-10 = -1.0460775e+18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101111100011101101100101000;
		b = 32'b11100011101100000110010000001101;
		correct = 32'b11101010001001101010010100110001;
		#400 //7739.3945 * -6.507673e+21 = -5.0365445e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011111110010011010001101010;
		b = 32'b10011100011101100000011101001000;
		correct = 32'b01010000111011110111111101110100;
		#400 //-3.9488068e+31 * -8.1403983e-22 = 32144860000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100111000000000010001011100;
		b = 32'b01111010101001111110111000010110;
		correct = 32'b11100000000100101111001100101111;
		#400 //-9.71519e-17 * 4.3597127e+35 = -4.2355435e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101110011001000001000101100;
		b = 32'b11010011110000111101011011010100;
		correct = 32'b01111010000111000111001011000110;
		#400 //-1.207205e+23 * -1682245700000.0 = 2.0308155e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001001110101001010110011111;
		b = 32'b10101100111100001001111010011111;
		correct = 32'b10010110101011110101111111100001;
		#400 //4.1430072e-14 * -6.8388207e-12 = -2.8333283e-25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000010011111000010100010000;
		b = 32'b01110000111111001101110111100101;
		correct = 32'b01100001110011001111101011011011;
		#400 //7.5495254e-10 * 6.260678e+29 = 4.7265148e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110101111010011011001000101;
		b = 32'b10101100000010111100001110110111;
		correct = 32'b10110011010011101001101000111110;
		#400 //24219.135 * -1.9861732e-12 = -4.8103395e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110000010001011111110001110;
		b = 32'b11100011001111010100101100010000;
		correct = 32'b00111001110010100011101100001001;
		#400 //-1.1046437e-25 * -3.4918435e+21 = 0.00038572427
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110111010100011101101111110;
		b = 32'b00001010001000011000110100111100;
		correct = 32'b10011001100100111101000010100100;
		#400 //-1964883700.0 * 7.778431e-33 = -1.5283713e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110010010101100001001011110;
		b = 32'b11110110010001011100110000010011;
		correct = 32'b01000101000111001010100100110100;
		#400 //-2.4992007e-30 * -1.0029508e+33 = 2506.5752
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101000011010100001000101100;
		b = 32'b01111110111010001111111000000111;
		correct = 32'b11010100100000001001000000100011;
		#400 //-2.8526924e-26 * 1.5484994e+38 = -4417392000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011110011010010000110101101;
		b = 32'b10100111001110111011000111001101;
		correct = 32'b01000011100101100110011000010010;
		#400 //-1.1547879e+17 * -2.604785e-15 = 300.79742
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100010000111101111000001010;
		b = 32'b11001000101011011011100111011100;
		correct = 32'b00010101100001001110101101000001;
		#400 //-1.5089071e-31 * -355790.88 = 5.368554e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001011010011000111000010000;
		b = 32'b10001001111001010111011111001111;
		correct = 32'b00111011110100010101100101100010;
		#400 //-1.156508e+30 * -5.5242412e-33 = 0.006388829
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100100110010110000010101111;
		b = 32'b00100110000100000100010000000000;
		correct = 32'b11011011001011001101111001000000;
		#400 //-9.721465e+31 * 5.0052193e-16 = -4.8658062e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000110000110000000111010101;
		b = 32'b01111001000110110011001110101011;
		correct = 32'b01000010011011000111001011101111;
		#400 //1.1736566e-33 * 5.0365873e+34 = 59.11224
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000100110110101110010101100;
		b = 32'b00101101001010110010000010001101;
		correct = 32'b00000110010011111011010101010000;
		#400 //4.0160136e-24 * 9.727452e-12 = 3.906558e-35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001000001011110100101001010;
		b = 32'b10110101110001111111001001111000;
		correct = 32'b01011111010100010010111001011100;
		#400 //-1.0118051e+25 * -1.4897223e-06 = 1.5073086e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001100010011111101011101101;
		b = 32'b10000111110110010010001100010000;
		correct = 32'b01000001111010100001000100110010;
		#400 //-8.955426e+34 * -3.267114e-34 = 29.258396
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001111010110010111010101100;
		b = 32'b01001101001110101011001001101101;
		correct = 32'b00001111101010111000001111010100;
		#400 //8.639234e-38 * 195765970.0 = 1.691268e-29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111010000000001111010001000;
		b = 32'b00000011011100110101110011100011;
		correct = 32'b10111011001101101010001010110000;
		#400 //-3.8966416e+33 * 7.151791e-37 = -0.0027867965
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001110001110000011101100110;
		b = 32'b01001111001100100010011100001101;
		correct = 32'b01010001100010101000000110000001;
		#400 //24.878613 * 2988903700.0 = 74359775000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101110101111100001100010101;
		b = 32'b00011101011011111000101001111000;
		correct = 32'b00101011110010011110001111010101;
		#400 //452485800.0 * 3.1702973e-21 = 1.4345145e-12
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101110101101000001111010110;
		b = 32'b10100101011111110000000011011011;
		correct = 32'b01011011110101011010111000001010;
		#400 //-5.438601e+32 * -2.2118014e-16 = 1.2029106e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000000101100111010110011111;
		b = 32'b01000110001101110110000101001100;
		correct = 32'b10011110110101111000111010001000;
		#400 //-1.944643e-24 * 11736.324 = -2.282296e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101011001100111101110110101;
		b = 32'b00010011010001010111000110001111;
		correct = 32'b00011001001100011100001101110000;
		#400 //3687.7317 * 2.4920884e-27 = 9.190154e-24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011110111001111111101001001;
		b = 32'b11100010111010101010000110100000;
		correct = 32'b10110111010010101000110011011111;
		#400 //5.578754e-27 * -2.1640922e+21 = -1.2072937e-05
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111100011110101100011110001;
		b = 32'b10101101001100101010101110100010;
		correct = 32'b00101101010010000001011111100101;
		#400 //-1.1199018 * -1.0156239e-11 = 1.1373989e-11
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010110110000111101011001110;
		b = 32'b11101000010100101000011110100011;
		correct = 32'b01110011101100100000011101110000;
		#400 //-7093607.0 * -3.976796e+24 = 2.820983e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101000110010101110101111101;
		b = 32'b11100011000101110001000001101001;
		correct = 32'b11100000101101001111111111110011;
		#400 //0.037442673 * -2.7866408e+21 = -1.0433928e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111000001000111011111110100111;
		b = 32'b00111100100000100000110001000110;
		correct = 32'b00110101001001100101111001011001;
		#400 //3.904072e-05 * 0.015874993 = 6.1977113e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101110011111110110000011111;
		b = 32'b01100111000000011000100100110111;
		correct = 32'b01100101010100100110101011011011;
		#400 //0.101524584 * 6.1171644e+23 = 6.2104256e+22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110110010011101011100101000;
		b = 32'b01000100100111001001011011010110;
		correct = 32'b00110011111101101110110000010010;
		#400 //9.178641e-11 * 1252.7136 = 1.14982086e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111100100100010101101011110;
		b = 32'b01010011000100011010110001111000;
		correct = 32'b11101011001001100101101000010100;
		#400 //-321429900000000.0 * 625663800000.0 = -2.0110707e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100011110010010111010011100;
		b = 32'b10000101101110100001000011011111;
		correct = 32'b00010010101101010001110001001001;
		#400 //-65321584.0 * -1.7497553e-35 = 1.1429679e-27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000001110100111110011111100;
		b = 32'b11000001111101111100101010010000;
		correct = 32'b11101010101101001000001000100111;
		#400 //3.522663e+24 * -30.973907 = -1.0911064e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011000011011010111000110001;
		b = 32'b11010010110110101011101011000100;
		correct = 32'b01011110011100100001101101100110;
		#400 //-9285169.0 * -469718140000.0 = 4.3614124e+18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000110100111100100110001001;
		b = 32'b00110000111010100101111000111000;
		correct = 32'b00011010010000011110010000101010;
		#400 //2.3513108e-14 * 1.7052519e-09 = 4.0095774e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110110101010100011000000101;
		b = 32'b01101010110100101011110111110000;
		correct = 32'b11100010001011111001000110101101;
		#400 //-6.356046e-06 * 1.2738569e+26 = -8.096693e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101100111101110100101101000;
		b = 32'b10100111001110001101110000000001;
		correct = 32'b11001101011001011000000010101000;
		#400 //9.380494e+22 * -2.5654394e-15 = -240650880.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011001001001001011000010101;
		b = 32'b10110001010011010111100011011010;
		correct = 32'b11000101000001000001100111100001;
		#400 //706892600000.0 * -2.9900122e-09 = -2113.6174
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000010111110010100111110110;
		b = 32'b11000110111101001011011001111000;
		correct = 32'b10110111110101010101001100001111;
		#400 //8.118656e-10 * -31323.234 = -2.5430256e-05
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100010110100011011100001111;
		b = 32'b11000011000100001011100100111100;
		correct = 32'b01101111111101101011100110111011;
		#400 //-1.05522334e+27 * -144.72357 = 1.5271569e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100100010111010011010011110;
		b = 32'b01101110010111101010100011101001;
		correct = 32'b11001011011100101110110101000011;
		#400 //-9.241318e-22 * 1.7227468e+28 = -15920451.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111111010010110110011111110;
		b = 32'b01100001101010101101011000100101;
		correct = 32'b11000010000110111100010110100100;
		#400 //-9.885965e-20 * 3.9392215e+20 = -38.94301
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010000101010000101011101001;
		b = 32'b11101111101111011001001001000000;
		correct = 32'b01011010010111001011110001100111;
		#400 //-1.3237644e-13 * -1.1733894e+29 = 1.5532911e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000100110110101000011100011;
		b = 32'b01001000001101101111000001001111;
		correct = 32'b00101001010111011111101010011010;
		#400 //2.6311548e-19 * 187329.23 = 4.928922e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101101100000110100000011011;
		b = 32'b10111101100101100101111011110111;
		correct = 32'b01010011110011110011110011100001;
		#400 //-24245147000000.0 * -0.07342332 = 1780159200000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010011101001011001111101001;
		b = 32'b00100110010011100100010101111011;
		correct = 32'b10110001010001010010101100110000;
		#400 //-4009210.2 * 7.156477e-16 = -2.8691822e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110011111101001010100000110;
		b = 32'b11000111000111000011011100011000;
		correct = 32'b01010110000110110101100110011010;
		#400 //-1067794800.0 * -39991.094 = 42702285000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011100000100001110101111010;
		b = 32'b11111100000110111100011111001111;
		correct = 32'b01010000000111100101101011001110;
		#400 //-3.284568e-27 * -3.2354345e+36 = 10627004000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000111010011011101000000000;
		b = 32'b01010000011011101001101001100111;
		correct = 32'b10100001110110011101011111100100;
		#400 //-9.2188874e-29 * 16012385000.0 = -1.4761638e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110011000111000110011111111;
		b = 32'b10011011110101110110111111100000;
		correct = 32'b10110010101111110111111011011011;
		#400 //62548680000000.0 * -3.5641064e-22 = -2.2293014e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111011010110111000001010111;
		b = 32'b01111010010111100110000110110010;
		correct = 32'b11001010010011001000010101000101;
		#400 //-1.16080304e-29 * 2.8866785e+35 = -3350865.2
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101101111000100101110001001;
		b = 32'b10000110100010010100001000011101;
		correct = 32'b10001100110010011110101000011010;
		#400 //6025.442 * -5.1630817e-35 = -3.1109848e-31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110010110100011011101101100;
		b = 32'b10100101010100001111001010100110;
		correct = 32'b10111100001100100001101111011110;
		#400 //59982892000000.0 * -1.8123337e-16 = -0.010870902
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110001100101010110010101010;
		b = 32'b11011110011101000000001110100111;
		correct = 32'b01001101001010100100111100011111;
		#400 //-4.062587e-11 * -4.3957702e+18 = 178582000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001111011100001110001001010;
		b = 32'b00111011100101001100101010001111;
		correct = 32'b01101110000010100110010011000010;
		#400 //2.3581322e+30 * 0.0045407484 = 1.0707685e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100001011110000001100011111;
		b = 32'b01011011010010111111110110000100;
		correct = 32'b10101000000010110111010011001010;
		#400 //-1.3482449e-31 * 5.7418164e+16 = -7.741375e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100100111110010010001111100;
		b = 32'b10111101100001101001110110000101;
		correct = 32'b00111010101001110101111000001010;
		#400 //-0.019426577 * -0.06573013 = 0.0012769115
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101000000100011001101010101;
		b = 32'b11100000110011100011000010110010;
		correct = 32'b01101110010100011011110000100101;
		#400 //-136525140.0 * -1.1886057e+20 = 1.6227455e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110010110111000111100111001;
		b = 32'b00100101001011011110111101011001;
		correct = 32'b10111100000101010010110100010001;
		#400 //-60352046000000.0 * 1.5086452e-16 = -0.009104983
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000111001110011110110001001;
		b = 32'b01011110100000011010101100100110;
		correct = 32'b01101111111010100100000100110101;
		#400 //31036557000.0 * 4.671802e+18 = 1.4499665e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000001110110111100000010110;
		b = 32'b11010011111100001100111110010101;
		correct = 32'b01011100101100000101100010011000;
		#400 //-191968.34 * -2068549600000.0 = 3.9709605e+17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000100010011010101101011011;
		b = 32'b00111010100001111111100000101100;
		correct = 32'b00001011100100100011110110100101;
		#400 //5.4300987e-29 * 0.0010373644 = 5.6329907e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100100010011001010111101110;
		b = 32'b11100110000010100111011111010111;
		correct = 32'b01101011000101001101011001110101;
		#400 //-1100.6853 * -1.634743e+23 = 1.7993377e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011110111101010110000110011;
		b = 32'b11010100011001000100000111000101;
		correct = 32'b01100000110001101000101010010010;
		#400 //-29186150.0 * -3921424000000.0 = 1.1445126e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100101000000000001010010000;
		b = 32'b00100110001011011111001100111110;
		correct = 32'b10111011010110010111001110001001;
		#400 //-5497902000000.0 * 6.0351087e-16 = -0.0033180437
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101000100111100110101000000;
		b = 32'b00101100111110001101000000111101;
		correct = 32'b00000010100011111010011100010000;
		#400 //2.9848327e-26 * 7.071703e-12 = 2.110785e-37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100101111111100110000011001;
		b = 32'b10101011100101000101000110100010;
		correct = 32'b00010000110111100011111001001111;
		#400 //-8.31788e-17 * -1.053869e-12 = 8.765956e-29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110011010110001001010000100;
		b = 32'b01110000000001000011100100001000;
		correct = 32'b01101110111100101101001111010101;
		#400 //0.22956282 * 1.6368387e+29 = 3.757573e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010010001110010101110101111;
		b = 32'b00010110100100111101011101001001;
		correct = 32'b10100001011001100000101100101000;
		#400 //-3263211.8 * 2.3884995e-25 = -7.7941796e-19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000101101011001100000010000;
		b = 32'b10100100111100111100001100101101;
		correct = 32'b10000110001011001110100111001010;
		#400 //3.076322e-19 * -1.0571509e-16 = -3.2521366e-35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011000010100110100010101110;
		b = 32'b00100110010001010000101010001100;
		correct = 32'b10110001110101010001000010000011;
		#400 //-9070766.0 * 6.83624e-16 = -6.200993e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001101010011001100110110100100;
		b = 32'b00111010011010110001100001101000;
		correct = 32'b00001000001111000001010001001100;
		#400 //6.3109884e-31 * 0.00089681754 = 5.659805e-34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101110001101101111011101111;
		b = 32'b11011001011111100000111000100010;
		correct = 32'b11010111110001010101110000101100;
		#400 //0.0971049 * -4469386500000000.0 = -433999330000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101101011010010001101101001;
		b = 32'b10011000000110001000101100101110;
		correct = 32'b10100110010011100101011001001111;
		#400 //363097380.0 * -1.9715807e-24 = -7.1587577e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011000010010110100101111000;
		b = 32'b11001011110000011011010100011001;
		correct = 32'b01010111010011111111001101110001;
		#400 //-9005432.0 * -25389618.0 = 228644480000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101001011100101000100000100;
		b = 32'b10011001111010100111001001100011;
		correct = 32'b00110111100111111010001111110001;
		#400 //-7.850516e+17 * -2.4241233e-23 = 1.9030618e-05
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110111101111101001000011101;
		b = 32'b10101100110100001011000100001111;
		correct = 32'b11000100010010100000011000011110;
		#400 //136240900000000.0 * -5.931373e-12 = -808.0956
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111010001000100001100100110;
		b = 32'b11000101110011010010001001111000;
		correct = 32'b00110101100111010100010000110010;
		#400 //-1.7849952e-10 * -6564.3086 = 1.1717259e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110010000010001111111010011;
		b = 32'b00111011100001101000101110011010;
		correct = 32'b00101010010010101111111111110010;
		#400 //4.3911385e-11 * 0.0041059973 = 1.8030003e-13
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110110100001011001001110100;
		b = 32'b10010101111101011101110100101111;
		correct = 32'b10010101010010000110111100011001;
		#400 //0.4076115 * -9.930368e-26 = -4.047732e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000011100110110010100010110;
		b = 32'b00111111111000100100011110101110;
		correct = 32'b10111000110101110010001101100100;
		#400 //-5.802986e-05 * 1.7678125 = -0.00010258591
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100010111010100001111100011;
		b = 32'b01010110100110100100001111101101;
		correct = 32'b11100011100001010101010110001100;
		#400 //-58003340.0 * 84808265000000.0 = -4.9191625e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000101001011100100100111000;
		b = 32'b00010000100111110000010110011000;
		correct = 32'b00010001110011011111011100110010;
		#400 //5.180813 * 6.272306e-29 = 3.2495643e-28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101011000000101011010111000;
		b = 32'b00101000100100001111000111110001;
		correct = 32'b11100110011111100000100110011001;
		#400 //-1.8637334e+37 * 1.6092137e-14 = -2.9991453e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010010000110110010010101111;
		b = 32'b00001110010110011000000000010000;
		correct = 32'b10001001001001100000001000010111;
		#400 //-0.00074536627 * 2.6808975e-30 = -1.9982506e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000111001110111011000011001111;
		b = 32'b11010101000101001111101110011101;
		correct = 32'b00011100110110100111010101100010;
		#400 //-1.4120276e-34 * -10238024000000.0 = 1.4456373e-21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111000101011001110100101011;
		b = 32'b01100001101001000000010111001111;
		correct = 32'b11000001001111111011100000101001;
		#400 //-3.1681984e-20 * 3.7821057e+20 = -11.982461
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001100101100011110101101000;
		b = 32'b10011101000001101100110101011011;
		correct = 32'b00011111000111100011100101010010;
		#400 //-18.779984 * -1.7840919e-21 = 3.3505216e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110110110111001010110010001;
		b = 32'b11001000010000011101001011100111;
		correct = 32'b01101111101001100100000010101001;
		#400 //-5.1847864e+23 * -198475.61 = 1.0290536e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010101001110011000101101111;
		b = 32'b10111000101111001001100011011000;
		correct = 32'b00100011111101100101100001000000;
		#400 //-2.969946e-13 * -8.993008e-05 = 2.6708749e-17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000110010010000001101100010;
		b = 32'b11011110010010110010011111010110;
		correct = 32'b01101111100111111000010011110110;
		#400 //-26979537000.0 * -3.659726e+18 = 9.873771e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011011000011110101001001111;
		b = 32'b11111100011001011100001100100000;
		correct = 32'b01000000010010101100001011001010;
		#400 //-6.639053e-37 * -4.7719743e+36 = 3.168139
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001000110001111101101000101;
		b = 32'b10101100001101010101000011100000;
		correct = 32'b11100101110110001011001111111000;
		#400 //4.964534e+34 * -2.5766542e-12 = -1.27918875e+23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101111010010001001101101110;
		b = 32'b10001001011110011100001010100000;
		correct = 32'b10010111111000110110010100011000;
		#400 //488795600.0 * -3.0063797e-33 = -1.4695051e-24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010101100000001111110000000;
		b = 32'b11101001100101110100011110110110;
		correct = 32'b11111100110100000010011111010101;
		#400 //378221360000.0 * -2.2860806e+25 = -8.646445e+36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111000000111000011110111111;
		b = 32'b01010001110111111101101010001011;
		correct = 32'b10101001011001100000011100010001;
		#400 //-4.249972e-25 * 120180530000.0 = -5.1076388e-14
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011101111010111000111000110;
		b = 32'b01001010001100100011111100011010;
		correct = 32'b10100110100000111110011111001110;
		#400 //-3.1340952e-22 * 2920390.5 = -9.152782e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010010101111111011101111110;
		b = 32'b10010110011100110111111111111010;
		correct = 32'b10001001010011010110101111100011;
		#400 //1.257092e-08 * -1.9669766e-25 = -2.4726706e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100011110111000011011100111;
		b = 32'b11001010001110000101110111111011;
		correct = 32'b01000111001101010010010101001101;
		#400 //-0.015351987 * -3020670.8 = 46373.3
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111001110111000111001111111;
		b = 32'b00111101111001001101011011111011;
		correct = 32'b10001101101001111010100001101010;
		#400 //-9.2472556e-30 * 0.11173817 = -1.0332714e-30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101010111001111101110111100;
		b = 32'b10001100110110010001110000100001;
		correct = 32'b00100010101110110110100110101010;
		#400 //-15185859000000.0 * -3.3451073e-31 = 5.0798328e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000000001011100100111010111;
		b = 32'b01100111010110110100110101110101;
		correct = 32'b11011111111001010011100001001100;
		#400 //-3.189765e-05 * 1.0356271e+24 = -3.303407e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011011000110000001010000011;
		b = 32'b10010110111000010100101000000111;
		correct = 32'b10011010110001111100011011011010;
		#400 //227.00981 * -3.6397428e-25 = -8.262573e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001000000100101010011000100;
		b = 32'b11001001001100010010001010110010;
		correct = 32'b01101010101101000101110010001011;
		#400 //-1.5026155e+20 * -725547.1 = 1.09021835e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101100100101001000100101101;
		b = 32'b10010100110011111000000011101011;
		correct = 32'b10001010111011011001101001100101;
		#400 //1.0920099e-06 * -2.0952508e-26 = -2.2880347e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001111000101111100111011110;
		b = 32'b01000000011100010000101101101011;
		correct = 32'b01010010110101011011011101011010;
		#400 //121856836000.0 * 3.766322 = 458952080000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011001010000011110011111100;
		b = 32'b00010011001001110001011110011000;
		correct = 32'b11001110110110111001111010010100;
		#400 //-8.735428e+35 * 2.1089996e-27 = -1842301400.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111001000111110111101000111;
		b = 32'b10111001011110110011000011001111;
		correct = 32'b00010001001000001101101011011100;
		#400 //-5.297015e-25 * -0.00023955408 = 1.2689216e-28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010010011101101110101100000;
		b = 32'b00010001001001011000010100111100;
		correct = 32'b10101100000001011100000001011000;
		#400 //-1.4556812e+16 * 1.3057261e-28 = -1.900721e-12
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111010010101011011000001000;
		b = 32'b10111111010010000100100101110011;
		correct = 32'b10000111000111101001100001011111;
		#400 //1.5250285e-34 * -0.78237075 = -1.1931377e-34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110110010001011101101111010;
		b = 32'b00001100011001010000110110000011;
		correct = 32'b11001011101100111001101001001100;
		#400 //-1.3340952e+38 * 1.7645584e-31 = -23540888.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010110011000100101100101100;
		b = 32'b10110110100110000001101110100011;
		correct = 32'b00111001111100101100010101100000;
		#400 //-102.14682 * -4.5331703e-06 = 0.00046304893
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101000010001010111000011110;
		b = 32'b00110100110111110101000111001111;
		correct = 32'b01001010011011100111011010110011;
		#400 //9392588000000.0 * 4.159651e-07 = 3906988.8
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101001101111001111101110100;
		b = 32'b00100010101000111110000100000001;
		correct = 32'b01011000011010110001011111010101;
		#400 //2.3276963e+32 * 4.441947e-18 = 1033950360000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001100110000000100110110101;
		b = 32'b00111010101110111011101000010001;
		correct = 32'b01101100110111101111101100110001;
		#400 //1.5057106e+30 * 0.001432242 = 2.156542e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000010110110101001110010110;
		b = 32'b01100011000010001100010001111001;
		correct = 32'b01010011111010100101100101110111;
		#400 //7.979052e-10 * 2.5229145e+21 = 2013046600000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000010000011011100100111100;
		b = 32'b10100110110011111001101000110110;
		correct = 32'b11010111100111010001100101111010;
		#400 //2.3981817e+29 * -1.4405309e-15 = -345465500000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011011101111110001101000100;
		b = 32'b11001010010111101001001101010010;
		correct = 32'b11001110010101111000010110111100;
		#400 //247.88776 * -3646676.5 = -903966460.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110100110111101110000010100;
		b = 32'b01100110110010000101111010100100;
		correct = 32'b10111101111100111111101100011101;
		#400 //-2.518049e-25 * 4.7310955e+23 = -0.119131304
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010101110001010000011001110;
		b = 32'b00111111101111110000101101100101;
		correct = 32'b00100011000010011100100000110001;
		#400 //5.004356e-18 * 1.4925352 = 7.469177e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111011110100010011110001010;
		b = 32'b11101010111111110110001011100101;
		correct = 32'b01111010111110011000111000000101;
		#400 //-4196895200.0 * -1.5437155e+26 = 6.478812e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000100101010100000001100001010;
		b = 32'b01001001010001101000111111000110;
		correct = 32'b10001110100000111101110111010101;
		#400 //-3.99696e-36 * 813308.4 = -3.250761e-30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001100101110110000001110110;
		b = 32'b10101000101000111010111011111001;
		correct = 32'b01010010110000011001001111000100;
		#400 //-2.2875415e+25 * -1.8172518e-14 = 415703900000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001111100001101001011101001;
		b = 32'b01100111011101010001011110001000;
		correct = 32'b01100001111001101000111111111100;
		#400 //0.00045933507 * 1.15741386e+24 = 5.316408e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100100011001011011000111010;
		b = 32'b11111101101000100011100000110010;
		correct = 32'b11000010101100100101010001101000;
		#400 //3.308119e-36 * -2.695334e+37 = -89.164856
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000110000010011001111011001;
		b = 32'b00101000110100000010000100101110;
		correct = 32'b11010010000111010001001100101011;
		#400 //-7.298985e+24 * 2.3107028e-14 = -168657860000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100001111111101011011010100;
		b = 32'b00101000010110111000111111011011;
		correct = 32'b11010101001001001000100010010100;
		#400 //-9.276773e+26 * 1.2188136e-14 = -11306657000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000001000001010101111001011;
		b = 32'b01010111000000000011111101011001;
		correct = 32'b01011111101000001111101101001111;
		#400 //164527.17 * 141009560000000.0 = 2.3199904e+19
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101111101100101010101000010;
		b = 32'b11001001000000010001111110001110;
		correct = 32'b11110111011110000111111010100110;
		#400 //9.529548e+27 * -528888.9 = -5.0400717e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001111110110111100010101100;
		b = 32'b01011001010000110100110011111011;
		correct = 32'b01110011101111111101100010001001;
		#400 //8847862400000000.0 * 3435766300000000.0 = 3.0399187e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101011101111010111001011001;
		b = 32'b11110011100001101110111101111000;
		correct = 32'b11101001100000101000110011110010;
		#400 //9.226838e-07 * -2.1381372e+31 = -1.9728244e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010011101000010101110000101;
		b = 32'b01000101101001001010011001101100;
		correct = 32'b01111000100111010000101010011100;
		#400 //4.836285e+30 * 5268.8027 = 2.548143e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101100010111101010011111111;
		b = 32'b00011010011111011101001000100011;
		correct = 32'b10011000100010101010010001001000;
		#400 //-0.06827735 * 5.248892e-23 = -3.5838046e-24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111111010101000010100000010;
		b = 32'b11001000011001011101010011011101;
		correct = 32'b11000000110100101000101111111011;
		#400 //2.795691e-05 * -235347.45 = -6.5795875
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110111001110110100001111001;
		b = 32'b00010110111011100000110100101001;
		correct = 32'b11001110010101110010111100000110;
		#400 //-2.3467569e+33 * 3.845928e-25 = -902545800.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010111110001100010101001101;
		b = 32'b11111110110001011011100111011100;
		correct = 32'b01011010010000000010010001110001;
		#400 //-1.0288915e-22 * -1.3141148e+38 = 1.3520816e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001010101011010111000000000;
		b = 32'b01011010111000100100011001101101;
		correct = 32'b11001100101111001101111001100101;
		#400 //-3.1094487e-09 * 3.184539e+16 = -99021610.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001011000111000101001010000;
		b = 32'b10010110110011001001010111101110;
		correct = 32'b10000000101101011101011101111011;
		#400 //5.0524092e-14 * -3.3052596e-25 = -1.6699525e-38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001110110110010011010101110;
		b = 32'b01010111011000110101100101110101;
		correct = 32'b11101001110000101001111111100001;
		#400 //-117655850000.0 * 249973350000000.0 = -2.9410827e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110110000011011110110000010;
		b = 32'b11001110000110010010010010111010;
		correct = 32'b00011101011001111100110000011100;
		#400 //-4.7760663e-30 * -642330240.0 = 3.0678118e-21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000010010100101010011101100;
		b = 32'b10111100110001101010001010110100;
		correct = 32'b10001101100111001111111001000111;
		#400 //3.9902897e-29 * -0.024247505 = -9.675457e-31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001101101101011100001111011;
		b = 32'b11101000000111010001000111111100;
		correct = 32'b01111010011000000011011111110011;
		#400 //-98097390000.0 * -2.9669732e+24 = 2.9105232e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010001111110101100100100010;
		b = 32'b01010100110010001100011010000101;
		correct = 32'b11010111100101100001001000000101;
		#400 //-47.837044 * 6898592500000.0 = -330008270000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111110011111001001011010101;
		b = 32'b10011011001000001101011011110010;
		correct = 32'b00100011100000100110101000001110;
		#400 //-106277.664 * -1.3304342e-22 = 1.4139544e-17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100011100011011011011001100;
		b = 32'b01010000111010000000101000110011;
		correct = 32'b00011101110110110001011101001010;
		#400 //1.8620973e-31 * 31143860000.0 = 5.7992898e-21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001001010101100101110001101;
		b = 32'b11001110111111000011010010111000;
		correct = 32'b10011000101010000100001110001011;
		#400 //2.0558715e-33 * -2115656700.0 = -4.3495183e-24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010110111001001110111010000;
		b = 32'b01010111011110000001101011000000;
		correct = 32'b11000010110101011100111111101111;
		#400 //-3.9189355e-13 * 272793770000000.0 = -106.90612
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110001010011110001011100110;
		b = 32'b00101010010110010000110001101101;
		correct = 32'b01010001000100000000100110010100;
		#400 //2.0056637e+23 * 1.9277783e-13 = 38664750000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000001011000111111000100110;
		b = 32'b00011100001100010011000010001111;
		correct = 32'b10110100111011101100011111100001;
		#400 //-758631200000000.0 * 5.862715e-22 = -4.4476386e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011111110101010110101011000;
		b = 32'b00101101011000010101001111100011;
		correct = 32'b00001001110111001010010001111111;
		#400 //4.1471051e-22 * 1.2808396e-11 = 5.3117765e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001100101000100110010000110;
		b = 32'b00011111001110110000111001111001;
		correct = 32'b10000001010110001011100010010000;
		#400 //-1.0049126e-18 * 3.9610762e-20 = -3.9805351e-38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100100111110100000000010110;
		b = 32'b00100001001110001011101101011001;
		correct = 32'b01000110011001011101010100110110;
		#400 //2.3501201e+22 * 6.258958e-19 = 14709.303
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000111011011110100100010110101;
		b = 32'b01010100111001001111100110101010;
		correct = 32'b10011100110101100000011000011110;
		#400 //-1.8001728e-34 * 7867529700000.0 = -1.4162913e-21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011001110100100010101111000;
		b = 32'b01111010110111001011011101110010;
		correct = 32'b01110110101000001001100100101110;
		#400 //0.0028422754 * 5.73013e+35 = 1.6286608e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001010001100011100010000011;
		b = 32'b10100111101010110001111110101000;
		correct = 32'b11000001100001001000000001000010;
		#400 //3487136300000000.0 * -4.7496356e-15 = -16.562626
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101101110001000010001010010111;
		b = 32'b01100101111010101011000010100111;
		correct = 32'b01010100001100111100111011110110;
		#400 //2.2297981e-11 * 1.3853655e+23 = 3089085500000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101011011100101111000101101;
		b = 32'b00010000000101000010001101010000;
		correct = 32'b10011110000010011110111101010011;
		#400 //-249946830.0 * 2.9215057e-29 = -7.302211e-21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101111100010010011110110100;
		b = 32'b01100001110001101110001010000001;
		correct = 32'b11110000001110110101101000010100;
		#400 //-505738880.0 * 4.5859708e+20 = -2.3193038e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001101111101100011001101110;
		b = 32'b11011000100011101010110011110101;
		correct = 32'b11100010110101001010010111101010;
		#400 //1562829.8 * -1254988000000000.0 = -1.9613326e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011001100101000100000111111;
		b = 32'b10111101000011101011010011111101;
		correct = 32'b00001000110001110000101110010110;
		#400 //-3.4384053e-32 * -0.034840573 = 1.1979601e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101001100101011110000000010;
		b = 32'b01001001110101011100011100011111;
		correct = 32'b01101111100101010100000101110011;
		#400 //5.2753085e+22 * 1751267.9 = 9.238478e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111101000110001111011010000;
		b = 32'b10001101101011100000110011000001;
		correct = 32'b10000101110111011100111000100100;
		#400 //1.9445462e-05 * -1.0726648e-30 = -2.0858464e-35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100100011111001001111010010;
		b = 32'b00001100100011000011010110011110;
		correct = 32'b00001001100111010100010111010010;
		#400 //0.01752654 * 2.1602685e-31 = 3.7862034e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011001010101000100001100011;
		b = 32'b11011111001101100111000001010001;
		correct = 32'b00100010111100110000111110010000;
		#400 //-5.0115074e-37 * -1.3146096e+19 = 6.588176e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010111101111110010110011101;
		b = 32'b01011101100010001111101010101001;
		correct = 32'b01100001000001001010010010110101;
		#400 //123.94846 * 1.2337984e+18 = 1.5292741e+20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100001010001010111101100001;
		b = 32'b10111101100010010101110111010010;
		correct = 32'b01111010001101010000011101011010;
		#400 //-3.503452e+36 * -0.06707348 = 2.349887e+35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011001000110001001010111011;
		b = 32'b10101100101011000001101110111100;
		correct = 32'b11101000010110110100010010000001;
		#400 //8.467243e+35 * -4.891613e-12 = -4.1418477e+24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110101011111101001101001110;
		b = 32'b11101011000011001110100001100111;
		correct = 32'b01101010010000011000111001011010;
		#400 //-0.343409 * -1.703471e+26 = 5.849873e+25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001000100110100111001001100;
		b = 32'b01000101011100011110111001111111;
		correct = 32'b10101111000010110011010111110001;
		#400 //-3.270847e-14 * 3870.906 = -1.266114e-10
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101010100111000010101010000;
		b = 32'b00111101010100011010010010010001;
		correct = 32'b00110011001011010011011111010000;
		#400 //7.879762e-07 * 0.051182333 = 4.0330463e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000111011000010000100000111;
		b = 32'b10001010010000101110010010100111;
		correct = 32'b10001011101100111100001111101111;
		#400 //7.3790317 * -9.383765e-33 = -6.92431e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000010110010100010001000110;
		b = 32'b11011011100010110011011011000110;
		correct = 32'b10110100011011000100110100011101;
		#400 //2.8081062e-24 * -7.837049e+16 = -2.2007266e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010110100110000110011111011;
		b = 32'b11011100000001100011100000011010;
		correct = 32'b11100111010111010100111000010111;
		#400 //6915709.5 * -1.5111732e+17 = -1.0450835e+24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011100110011111110100111100;
		b = 32'b10010001000111101111101011100001;
		correct = 32'b00010101001111110100001001100111;
		#400 //-307.9784 * -1.254131e-28 = 3.8624525e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001110001010111101110101010;
		b = 32'b11000111111000100011000010001110;
		correct = 32'b10110010001011100111110010100001;
		#400 //8.77001e-14 * -115809.11 = -1.015647e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100001010111011011011011101;
		b = 32'b11000010011001101101010001110111;
		correct = 32'b11001111000110101101010011001110;
		#400 //45013876.0 * -57.707485 = -2597637600.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001010011001100011000011001;
		b = 32'b10000000110110001110101111100100;
		correct = 32'b10111010101011011000001111010101;
		#400 //6.6452904e+34 * -1.9921089e-38 = -0.0013238142
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110111111110100010010100101;
		b = 32'b01010110101110100001000101111001;
		correct = 32'b01010110001110011000100101001100;
		#400 //0.4985706 * 102292100000000.0 = 50999834000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011001110111000110101000101;
		b = 32'b01101000000100011000100011010111;
		correct = 32'b01010011110101010011111010001001;
		#400 //6.6631797e-13 * 2.7490696e+24 = 1831754400000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001000111100111010111111000;
		b = 32'b01100011100010101001010101110011;
		correct = 32'b01101101001010111001000000110011;
		#400 //649055.5 * 5.112839e+21 = 3.3185164e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011001010010111010000110111;
		b = 32'b01111011001101101110000110010000;
		correct = 32'b01101110111100100001101111011011;
		#400 //3.9454076e-08 * 9.49573e+35 = 3.7464524e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100011011101101011001010100;
		b = 32'b00111001111111000000100101100001;
		correct = 32'b10110110111010110010001110111011;
		#400 //-0.014577467 * 0.00048072173 = -7.0077053e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001100010110111111001100100;
		b = 32'b00010100111010100111000111111110;
		correct = 32'b10000110111111110111111101001001;
		#400 //-4.0598014e-09 * 2.3672924e-26 = -9.610737e-35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010110110101011110000001011;
		b = 32'b11001010001010001110000100111000;
		correct = 32'b00110101100100000100101111010110;
		#400 //-3.885506e-13 * -2766926.0 = 1.0750907e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000001110000111110001011011;
		b = 32'b01000100010101000011101000010001;
		correct = 32'b11101101000110001111000011010100;
		#400 //-3.4848375e+24 * 848.9073 = -2.958304e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000000100111101100101010001;
		b = 32'b10100011101101001010101001010010;
		correct = 32'b00000100010100001010111001010101;
		#400 //-1.2523288e-19 * -1.9587773e-17 = 2.4530332e-36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100001110010100111000000101;
		b = 32'b11111000010110111101110011001000;
		correct = 32'b01100101000111110010010110001110;
		#400 //-2.633339e-12 * -1.7837359e+34 = 4.6971815e+22
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111110000011100110001011111;
		b = 32'b00100101000101001111111011011110;
		correct = 32'b10100101011000011001011000110000;
		#400 //-1.5140494 * 1.2923306e-16 = -1.9566525e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010010100010101111100100110;
		b = 32'b00101000001101111011001001011010;
		correct = 32'b01001011000101100011110011100010;
		#400 //9.655564e+20 * 1.01972145e-14 = 9845986.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110001101001100110010110011;
		b = 32'b01011011101110110110111101111001;
		correct = 32'b11110010100001000110000001000001;
		#400 //-49697817000000.0 * 1.0551677e+17 = -5.243953e+30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111001100110100111001101100;
		b = 32'b10110001111101110010001000001000;
		correct = 32'b00010001101011010001100010000000;
		#400 //-3.7969593e-20 * -7.192515e-09 = 2.7309687e-28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110011011010110101000011000;
		b = 32'b01000101011011110110000011110011;
		correct = 32'b10111100010111011111111111110110;
		#400 //-3.5377507e-06 * 3830.0593 = -0.013549795
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110101101000110011111111000;
		b = 32'b10011110110011001000110110111111;
		correct = 32'b10100110000100000010011010111101;
		#400 //23091.984 * -2.1657965e-20 = -5.0012536e-16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011010101001010101000011000;
		b = 32'b00010010001110100000101111110110;
		correct = 32'b10111110000110101000110110000101;
		#400 //-2.5709552e+26 * 5.8705994e-28 = -0.15093048
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000111101111011111111000100;
		b = 32'b01110011011011110000000011010101;
		correct = 32'b11001100111001110100110011010110;
		#400 //-6.4041637e-24 * 1.8935788e+31 = -121267890.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010100100001110110111101011;
		b = 32'b00110110001001001010100100011100;
		correct = 32'b00110001001110100111000001001111;
		#400 //0.0011057233 * 2.453634e-06 = 2.7130402e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111101000000000110110110011;
		b = 32'b00011101111111101110110000110001;
		correct = 32'b01000110000111110110000101000011;
		#400 //1.5116627e+24 * 6.7477456e-21 = 10200.315
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011010101110101110010100010;
		b = 32'b01011101001100001101101001100110;
		correct = 32'b11110001000101001100011101101010;
		#400 //-924972100000.0 * 7.9647564e+17 = -7.367177e+29
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100001000010110110101010100;
		b = 32'b11000110001011000000000110011001;
		correct = 32'b01001010110110001110110011101101;
		#400 //-645.70825 * -11008.399 = 7108214.5
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101001100000100100111110111;
		b = 32'b01110101001001001011101001101100;
		correct = 32'b00111010111000101101111110000101;
		#400 //8.2890654e-36 * 2.0881781e+32 = 0.0017309046
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111101011010010110101010001;
		b = 32'b10011101111011110001100010000000;
		correct = 32'b00001110001000011011110111100001;
		#400 //-3.1500716e-10 * -6.3288106e-21 = 1.9936206e-30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111010110101010010110110011;
		b = 32'b00101110011000001010011010010110;
		correct = 32'b01101110001111111101111101000100;
		#400 //2.9063206e+38 * 5.107966e-11 = 1.4845387e+28
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100110100110110000101011100;
		b = 32'b11100000110010111000011000111010;
		correct = 32'b10111110001010000000110100001001;
		#400 //1.3987976e-21 * -1.1732378e+20 = -0.16411223
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011011011101101111011000110;
		b = 32'b00110010110010111000001001001111;
		correct = 32'b00101110101111011110010000111110;
		#400 //0.0036448701 * 2.3691568e-08 = 8.635269e-11
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000100001011000100110100010;
		b = 32'b11010010000000011011011101111001;
		correct = 32'b11010011000001110101010000011110;
		#400 //4.173051 * -139282240000.0 = -581231840000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100111010001101111111100101;
		b = 32'b10110101011100100011001000000010;
		correct = 32'b01100010110111000101000100100100;
		#400 //-2.2522248e+27 * -9.0224796e-07 = 2.0320652e+21
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001000101110011001011110101;
		b = 32'b11010010011001100100110101010110;
		correct = 32'b10010100000010000000010101110101;
		#400 //2.777088e-38 * -247284990000.0 = -6.8673215e-27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001000011100101111000100110;
		b = 32'b11011001100111111010111101000101;
		correct = 32'b01010011001100011001101111100101;
		#400 //-0.00013577248 * -5618404000000000.0 = 762824700000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110101110100100001101100100;
		b = 32'b01001011000110110011100001000101;
		correct = 32'b01010010011000011101111101111101;
		#400 //23841.695 * 10172485.0 = 242529290000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101111110100110001101111110;
		b = 32'b11011100111011110100100111111001;
		correct = 32'b00101011011010100000101100111101;
		#400 //-1.5431391e-30 * -5.3883083e+17 = 8.3149096e-13
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001110000001100110000111111;
		b = 32'b11011001101101011110100001011000;
		correct = 32'b10110100000010001111111101100100;
		#400 //1.9934829e-23 * -6400304400000000.0 = -1.2758898e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110101111110110100101000110;
		b = 32'b00101111011011000000110001111011;
		correct = 32'b00010110101100000111111001100001;
		#400 //1.3281822e-15 * 2.1468509e-10 = 2.851409e-25
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011101001000100111100011011;
		b = 32'b11111101000101110000001101111001;
		correct = 32'b01111001010000011101100111000111;
		#400 //-0.005014313 * -1.2545716e+37 = 6.2908146e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000111000111011010010101100;
		b = 32'b11011011000110101101100011101101;
		correct = 32'b00111100100010011011101110100011;
		#400 //-3.8574854e-19 * -4.358566e+16 = 0.016813105
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100111111010110010001001000;
		b = 32'b11001001010010110101110001011100;
		correct = 32'b10001110110010010100100111110000;
		#400 //5.9572108e-36 * -832965.75 = -4.9621525e-30
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010100110001010110010101010;
		b = 32'b10011011001011011011100110000111;
		correct = 32'b00011110010011110011011010101000;
		#400 //-76.337234 * -1.4370172e-22 = 1.0969791e-20
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111010001001110011101000000;
		b = 32'b01001100001100110001011011010101;
		correct = 32'b10110100000010011011111101000001;
		#400 //-2.7325825e-15 * 46947156.0 = -1.2828697e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001100111111110110011000100;
		b = 32'b11011000010001010110000000100010;
		correct = 32'b11010010011101101001101010000010;
		#400 //0.00030503247 * -868066700000000.0 = -264788540000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010110010000011110000100111;
		b = 32'b11010110011101110010001000111100;
		correct = 32'b00110001110000010100110011010001;
		#400 //-8.281524e-23 * -67931600000000.0 = 5.6257723e-09
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110110001111110101101101000100;
		b = 32'b00010101100101100001101011101001;
		correct = 32'b01001100011000000110011100101111;
		#400 //9.7029276e+32 * 6.0626974e-26 = 58825916.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100101110101101011110001101;
		b = 32'b10010010011101010011110000111000;
		correct = 32'b00111111101100101111110000111101;
		#400 //-1.8070249e+27 * -7.7382594e-28 = 1.3983227
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100111100101101001011100110;
		b = 32'b01100101111011011000000011000011;
		correct = 32'b01111011011000010100011101100001;
		#400 //8343363000000.0 * 1.4019701e+23 = 1.1697145e+36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001101110010011100000011001;
		b = 32'b11100111011100011101001100001110;
		correct = 32'b11010001101011101111011010000011;
		#400 //8.225382e-14 * -1.1419836e+24 = -93932510000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100001000100000011100000100;
		b = 32'b00000101110110000101100111101000;
		correct = 32'b10001010100010001110111011010011;
		#400 //-648.1096 * 2.0345569e-35 = -1.318616e-32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010110010011100011010101010;
		b = 32'b11100000011111010011101011000101;
		correct = 32'b10100011110001111001011110101000;
		#400 //2.9648323e-37 * -7.2988454e+19 = -2.1639852e-17
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111100000100000101010011000;
		b = 32'b11110000001011011011100000101011;
		correct = 32'b10111000001100000111110101101100;
		#400 //1.9566452e-34 * -2.150542e+29 = -4.2078478e-05
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111100010110100101111100010;
		b = 32'b10010010010100001101100111001010;
		correct = 32'b00100010011000110100100001010010;
		#400 //-4674012000.0 * -6.5901673e-28 = 3.0802523e-18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100011001010101001000110011;
		b = 32'b10001111010011111000101000111111;
		correct = 32'b10110100001110011110100101001110;
		#400 //1.692091e+22 * -1.0232513e-29 = -1.7314343e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110111101101000100001011101;
		b = 32'b01001000000100001100011001011111;
		correct = 32'b01100111100010110110101110111101;
		#400 //8.8822755e+18 * 148249.48 = 1.3167927e+24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111011010010011111001111000;
		b = 32'b10110110011110100000110001110111;
		correct = 32'b00111110011000111101001001011101;
		#400 //-59710.47 * -3.7260158e-06 = 0.22248216
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010101011111000101101011001;
		b = 32'b01000000111101011001001111100011;
		correct = 32'b01000100001010000110010111000101;
		#400 //87.77216 * 7.6743026 = 673.59015
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100111001010111010000000011;
		b = 32'b01011111000000101010110101110110;
		correct = 32'b10111100011010100100000011000101;
		#400 //-1.5183937e-21 * 9.416312e+18 = -0.014297669
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101110000101100001000001110;
		b = 32'b11110101010111001100010011011100;
		correct = 32'b11101011101001111111010010001000;
		#400 //1.4510604e-06 * -2.7985793e+32 = -4.0609076e+26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001000001011001000001000100;
		b = 32'b11101110000001001001111001111100;
		correct = 32'b01010111100010100110001000100110;
		#400 //-2.9657063e-14 * -1.0260904e+28 = 304308300000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000000101001010100101111001;
		b = 32'b11010100100011100011110010011101;
		correct = 32'b11110101001001010011001001101000;
		#400 //4.2848905e+19 * -4887218000000.0 = -2.0941195e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011001011001010110011101010;
		b = 32'b11110011010111001101110111110001;
		correct = 32'b01000111000101001111101001001101;
		#400 //-2.1794705e-27 * -1.7498883e+31 = 38138.3
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011000111100100101000001000;
		b = 32'b00111111101111001011111000001101;
		correct = 32'b01110011011010010110011111000010;
		#400 //1.2540961e+31 * 1.4745499 = 1.8492273e+31
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001010000010001000110101101;
		b = 32'b01110110110110110101010111111101;
		correct = 32'b01111000101001010110101011111001;
		#400 //12.066815 * 2.2243302e+33 = 2.6840583e+34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011010111011100110111110100;
		b = 32'b01000010011101101101110101101010;
		correct = 32'b00000110010101011110001110111111;
		#400 //6.5182485e-37 * 61.716225 = 4.022817e-35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010101001101101110000111111;
		b = 32'b11000011100010000010000111110101;
		correct = 32'b11110110101100010111011001000111;
		#400 //6.610019e+30 * -272.2653 = -1.7996787e+33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111000101011011010100011110;
		b = 32'b01101011001000010100111100110010;
		correct = 32'b11001010101111001010101001110000;
		#400 //-3.1701794e-20 * 1.9501105e+26 = -6182200.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110110110010011010010110110;
		b = 32'b11001010010000001010111111100010;
		correct = 32'b10011001101000110111110011000011;
		#400 //5.354539e-30 * -3156984.5 = -1.6904196e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010001100111110001011111101;
		b = 32'b11000010111111000111001100010011;
		correct = 32'b00010101101100010110010001001101;
		#400 //-5.6762225e-28 * -126.224754 = 7.164798e-26
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011100111101001101000011011;
		b = 32'b00011101010101110000101010110011;
		correct = 32'b00000001100001010011101000001110;
		#400 //1.719566e-17 * 2.8460544e-21 = 4.893979e-38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010111100111010111010011011;
		b = 32'b10111001010000101100010011110100;
		correct = 32'b01101100101110010110010111001011;
		#400 //-9.6532406e+30 * -0.00018574652 = 1.7930558e+27
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001011010000111101100000101;
		b = 32'b10001111100111111000101110001011;
		correct = 32'b10011001100100001110001100100001;
		#400 //952240.3 * -1.573236e-29 = -1.4980988e-23
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110000010110100110111001011;
		b = 32'b11011011100000111101101111011000;
		correct = 32'b00111010000011111000000011100000;
		#400 //-7.374686e-21 * -7.4229885e+16 = 0.0005474221
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010001010001010100001111011;
		b = 32'b00111101101000111001110101011010;
		correct = 32'b00001000010101111001010111100010;
		#400 //8.1205934e-33 * 0.07988997 = 6.4875395e-34
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011110010000100111101110010;
		b = 32'b10000111011101101110011000110000;
		correct = 32'b00111011110000010011000001110100;
		#400 //-3.174044e+31 * -1.8574629e-34 = 0.0058956686
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001011101011001001001100001;
		b = 32'b00100001011111011011011011100111;
		correct = 32'b00110011011100110110000100011110;
		#400 //65920176000.0 * 8.5961803e-19 = 5.6666174e-08
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000000100010001011100010001;
		b = 32'b01001000100010110110100011011111;
		correct = 32'b00111001000111100000010111101100;
		#400 //5.278347e-10 * 285510.97 = 0.0001507026
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011110110101100001010001010;
		b = 32'b10011011100011110110111000001000;
		correct = 32'b00100111111101010010000101100011;
		#400 //-28673300.0 * -2.3728472e-22 = 6.803736e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100011100000000000111100011;
		b = 32'b10100001011001000001010101000110;
		correct = 32'b01001110010101011101010110100000;
		#400 //-1.1606044e+27 * -7.727756e-19 = 896886800.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011101110001000100101101000;
		b = 32'b01010111000010000000011100011100;
		correct = 32'b11111011010001000001110000111110;
		#400 //-6.808204e+21 * 149564120000000.0 = -1.018263e+36
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111010100011100000100100100;
		b = 32'b00000000001000100101100000011011;
		correct = 32'b00100111011000010001111010111010;
		#400 //9.905374e+23 * 3.154013e-39 = 3.124168e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011110110111110110101110111;
		b = 32'b10100100110101011111100111001001;
		correct = 32'b11001001001101111101001100101011;
		#400 //8.113896e+21 * -9.279718e-17 = -752946.7
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010100000100000111110100101;
		b = 32'b11100101011010000001011000010101;
		correct = 32'b01011000011010111101001011001011;
		#400 //-1.5141106e-08 * -6.8499773e+22 = 1037162300000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101010001101111010001111111;
		b = 32'b01111101101001000010111100001010;
		correct = 32'b01011011011111110011001001100000;
		#400 //2.6331483e-21 * 2.7279704e+37 = 7.1831507e+16
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111100101110001100011111010;
		b = 32'b00010010000110001010101100011110;
		correct = 32'b10001010001101000011011110101000;
		#400 //-1.8012233e-05 * 4.817366e-28 = -8.6771525e-33
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000100001000111110000010001;
		b = 32'b01111100001100000001000110110001;
		correct = 32'b11110101001101100011110011100111;
		#400 //-6.31736e-05 * 3.6568123e+36 = -2.3101398e+32
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000000110111111110010001011;
		b = 32'b11101010011111110011010101001011;
		correct = 32'b01000011000110111000000100000111;
		#400 //-2.0160782e-24 * -7.713194e+25 = 155.50401
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101111001101101111101011010;
		b = 32'b10100000101011111111100001101000;
		correct = 32'b10101111000111101011001010110101;
		#400 //484174660.0 * -2.9810535e-19 = -1.4433506e-10
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011000010010101100010101001;
		b = 32'b10100011011010101101110011001101;
		correct = 32'b01001110111111000000001100000001;
		#400 //-1.6604152e+26 * -1.2731922e-17 = 2114027600.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011010000000110111011110101;
		b = 32'b11011010101101011000000111101101;
		correct = 32'b11010110100010000111000000011101;
		#400 //0.002936301 * -2.5544913e+16 = -75007550000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001001110110001010000100001;
		b = 32'b10010101001001001010110001010001;
		correct = 32'b10111110111100001010110110100100;
		#400 //1.4135262e+25 * -3.325547e-26 = -0.47007477
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011101101001000001100111111;
		b = 32'b00110000001010111010101010011100;
		correct = 32'b11010100011100100001011111110000;
		#400 //-6.6597424e+21 * 6.245189e-10 = -4159134800000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111110010111011101100010010;
		b = 32'b00110001100011110001101101101111;
		correct = 32'b00000001111000111100011010101000;
		#400 //2.0089402e-29 * 4.1649666e-09 = 8.367169e-38
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001110011001011001010100111;
		b = 32'b10011010101011111110001001011010;
		correct = 32'b11010101000011001010001100011110;
		#400 //1.3285651e+35 * -7.2743994e-23 = -9664513000000.0
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010100000001101011010101100;
		b = 32'b00010000100110001011000000101000;
		correct = 32'b10000011100110011011000000111100;
		#400 //-1.4998783e-08 * 6.022484e-29 = -9.032993e-37
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110000010010100111001001101;
		b = 32'b00110111100001100111000010110010;
		correct = 32'b11000110000100000011011011011100;
		#400 //-575902500.0 * 1.6026523e-05 = -9229.715
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010000111101001000100011111;
		b = 32'b00110011010001000111000010010111;
		correct = 32'b10000101111100110101100110110010;
		#400 //-5.0034885e-28 * 4.5737206e-08 = -2.2884559e-35
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101001001010111110010010001;
		b = 32'b10010001100010001110000011010010;
		correct = 32'b10100111001100001111011100000100;
		#400 //11372152000000.0 * -2.1595573e-28 = -2.4558814e-15
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010011010001001100111001001;
		b = 32'b00101011011011000010011100100001;
		correct = 32'b11000110010101101001000101010011;
		#400 //-1.6367821e+16 * 8.3898345e-13 = -13732.331
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000011110101110110011001101;
		b = 32'b00000110011111000110100001100101;
		correct = 32'b10110111011101110110011101101101;
		#400 //-3.106301e+29 * 4.747263e-35 = -1.4746428e-05
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001101010100010100001100100;
		b = 32'b11011011011111100000000100000111;
		correct = 32'b01011101101010001101010011000010;
		#400 //-21.269722 * -7.1495774e+16 = 1.5206952e+18
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101110011100111110001101111;
		b = 32'b00011001111100100011111110110110;
		correct = 32'b10011000010000110110010100000100;
		#400 //-0.100823276 * 2.5047946e-23 = -2.525416e-24
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010011111010001011100001000;
		b = 32'b01001001111110011011011110010100;
		correct = 32'b00110100111101101110000011100101;
		#400 //2.2478905e-13 * 2045682.5 = 4.5984703e-07
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100101001010010101000010001010;
		b = 32'b01001111111000110111100110001011;
		correct = 32'b10110101100101100111001011001101;
		#400 //-1.4685701e-16 * 7632787000.0 = -1.1209282e-06
					
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end

endmodule
