
    `include "alu.v"


    module or_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .A(a),
                .B(b),
                .OpCode(op),
                .O(out)
            );
        /* create a 10Mhz clock */
        always
        #100 clock = ~clock; // every 100 nanoseconds invert
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, a, b, op, out);
            clock = 0;

    op = 3'b101;

		/* Display the operation */
		$display ("Opcode: 101, Operation: OR");
		/* Test Cases!*/
		a = 32'b10100011101110110111010001110011;
		b = 32'b00101100010100101110001011011000;
		correct = 32'b10101111111110111111011011111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000101000001011100000101011;
		b = 32'b00000010100000111011001101101100;
		correct = 32'b11101010101000111011101101101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101101000100101101000001111;
		b = 32'b10101100011100001010010111001011;
		correct = 32'b10111101111100101111111111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010001100001000011110111011;
		b = 32'b01001111000100000110000011100101;
		correct = 32'b01111111001100001110011111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001100011110101100100010111;
		b = 32'b10011100010110011111101100111101;
		correct = 32'b11011101110111111111101100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001100010100110000110100111;
		b = 32'b00011111110101011000010110000010;
		correct = 32'b10111111110111111110010110100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110011101000011010000111000;
		b = 32'b11001011000100100110001001100000;
		correct = 32'b11001111011101100111011001111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110011010000100000101101110;
		b = 32'b11000000110110100111010000101101;
		correct = 32'b11100110111110100111010101101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100100000011100111111101111;
		b = 32'b01100001111100000110000010111111;
		correct = 32'b01110101111100011110111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100101011111100000110011111;
		b = 32'b00010111111100100100110100000010;
		correct = 32'b11110111111111111100110110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000000001110001010100001000;
		b = 32'b11011101001100000001101111010110;
		correct = 32'b11011101001101110001111111011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101000111000000010011001100;
		b = 32'b01001111100011001000000101000100;
		correct = 32'b11111111100111001000010111001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101000011100110000110001111;
		b = 32'b10000011100100001110010001110011;
		correct = 32'b10101111100111101110010111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100011011011111011010010000;
		b = 32'b10011011111100011110000101010100;
		correct = 32'b11011111111111011111011111010100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100111111100100111011110001;
		b = 32'b00010010100110100010010010010000;
		correct = 32'b10011110111111100110111011110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000101011101100001110010010;
		b = 32'b00000111101111100001010100000100;
		correct = 32'b10011111101111101101011110010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110000111000110000011011111;
		b = 32'b01101101100001011001101011001010;
		correct = 32'b11111111100111011111101011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111000000101110101111101110011;
		b = 32'b00111101001001111100101000101111;
		correct = 32'b11111101001101111101111101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101010000100100101011110101;
		b = 32'b01100001100000011101000000001011;
		correct = 32'b01100101110000111101101011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110100110111001001000101110;
		b = 32'b01100001100011101110000101111011;
		correct = 32'b01100111100111111111001101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001100001011011111001001010;
		b = 32'b00000010001110111011010011101001;
		correct = 32'b00100011101111111011111011101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011001010010111001100110010;
		b = 32'b11110011001000011110111000111110;
		correct = 32'b11110011001010011111111100111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110000111010010011110111101;
		b = 32'b10010000001000011001011100101010;
		correct = 32'b11111110001111011011011110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101110001011000001011110100;
		b = 32'b01111110010000110110111000010111;
		correct = 32'b01111111110001111110111011110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110001100010110101001111000;
		b = 32'b10111011110011100111010010001101;
		correct = 32'b10111111111111110111111011111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001000001100101101010111001;
		b = 32'b01111101111111000010000000110110;
		correct = 32'b01111101111111100111101010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111011101101111111011100000;
		b = 32'b11010010011111101010011101010101;
		correct = 32'b11011111011111101111111111110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010110010101101001111011100;
		b = 32'b11100111111111111101111101011001;
		correct = 32'b11100111111111111101111111011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101011111000001000000010001;
		b = 32'b10000101110011101010011111100111;
		correct = 32'b10011101111111101011011111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101100011011001110000011001;
		b = 32'b00100100000100001000110110101010;
		correct = 32'b11111101100111011001110110111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111000110000010110001100001110;
		b = 32'b10000100111100010111100110110101;
		correct = 32'b11111100111100010111101110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001110110011110000011110101;
		b = 32'b00010100011011111000101010100111;
		correct = 32'b10010101111111111110101011110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110000101100001001000010011;
		b = 32'b10110000100101010001100010000000;
		correct = 32'b11110110100101110001101010010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110001010010010000001001001;
		b = 32'b10010001101101011001001000000111;
		correct = 32'b11111111101111011011001001001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010000011111001000000011011;
		b = 32'b10110001100000000000110000110110;
		correct = 32'b10111011100011111001110000111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101100111101110110000000101;
		b = 32'b10010100010000110010101111000011;
		correct = 32'b11011101110111111110111111000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000011001100000100010111110;
		b = 32'b00110101000001111101011001001101;
		correct = 32'b01110101011001111101111011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110010101011001001101001001;
		b = 32'b01111110100111000011101001011010;
		correct = 32'b01111110110111011011101101011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111101010100010110110000100;
		b = 32'b01101001010101011010001011001111;
		correct = 32'b01101111111111111010111111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011011111000110101011011101;
		b = 32'b10100011111000111000111110001101;
		correct = 32'b11110011111111111110111111011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001111100100111110101000000;
		b = 32'b11110111000001001110110100001100;
		correct = 32'b11110111111101101111110101001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110001111000111000010011101;
		b = 32'b00011110101000010001010110110111;
		correct = 32'b00011110101111010111010110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000000000011110000101111010;
		b = 32'b10100101110001111101111011000110;
		correct = 32'b11111101110001111111111111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100011011011100010110000111;
		b = 32'b11101101000100100100110000010111;
		correct = 32'b11101101011111111100110110010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001010100110011100011111101;
		b = 32'b01011100000110000101111100001000;
		correct = 32'b11111101010110110111111111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010101101110011101100011000;
		b = 32'b00001001001111000100001110110000;
		correct = 32'b00111011101111110111101110111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010110010110010101011011101;
		b = 32'b11101011011011001111010110011110;
		correct = 32'b11101011111011111111111111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001111111000001000100010110;
		b = 32'b01111111001000011111100100111111;
		correct = 32'b01111111111111011111100100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011100111100111000100101110;
		b = 32'b00011111101110100110010101011101;
		correct = 32'b00011111101111100111010101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000111111100010110010101100;
		b = 32'b11100100110110001110110100000001;
		correct = 32'b11111100111111101110110110101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101000101101110101001101100;
		b = 32'b10101101101000010001101100101010;
		correct = 32'b10111101101101111111101101101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111111101100100000010011100;
		b = 32'b00100110110111001100110100000010;
		correct = 32'b10110111111111101100110110011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100010110101000100101001001;
		b = 32'b11111111110100111111000001101000;
		correct = 32'b11111111110110111111100101101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101110111011000000001010011;
		b = 32'b00000110110110010010100111100000;
		correct = 32'b01000111110111011010100111110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000110011100010111110011101;
		b = 32'b11111100000011111101100010000010;
		correct = 32'b11111100110011111111111110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111100000011110101010001111;
		b = 32'b10010101000010011000110010101010;
		correct = 32'b10010111100010011110111010101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101010111110001100100110000;
		b = 32'b00000101101111110000110010100011;
		correct = 32'b01110101111111110001110110110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100111110111110101011010101;
		b = 32'b10010100110010111100100111000111;
		correct = 32'b10111100111110111110101111010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001101111111011001010011101;
		b = 32'b10101000100111110101011010100100;
		correct = 32'b11101001101111111111011010111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010011010111000000101100110;
		b = 32'b10011101001001001100110010111100;
		correct = 32'b11011111011011111100110111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001100110111110011110100111;
		b = 32'b10100010101000011000010111110001;
		correct = 32'b11110011101110111110011111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000100001010100101000000011;
		b = 32'b11110011011110110011000110011110;
		correct = 32'b11111011111111110111101110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111101111000000111010110011;
		b = 32'b10000101111010110111111111000111;
		correct = 32'b11000111111111110111111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101101111111010101001110111011;
		b = 32'b11111000010100111111000111011010;
		correct = 32'b11111101111111111111001111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110000011011010111101111001;
		b = 32'b11101011101101100010011010000100;
		correct = 32'b11101111101111111010111111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001001010011111100100001001;
		b = 32'b10000010111000001000001011110001;
		correct = 32'b11000011111010011111101111111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110111010111010101100000000;
		b = 32'b10100010000011101110101001011000;
		correct = 32'b11100110111011111110101101011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101101101101101000000101011000;
		b = 32'b11001100110011011000000000101101;
		correct = 32'b11101101111111111000000101111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010011101111101010010100000;
		b = 32'b00011101100011001101111011100110;
		correct = 32'b11011111111111111101111011100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000101101110000000100000111;
		b = 32'b10100100101000100110111111001110;
		correct = 32'b10111100101101110110111111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000010111000011000110100111;
		b = 32'b10010111111101110011010001000010;
		correct = 32'b10011111111111110011010111100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010011010011110010100001101;
		b = 32'b00010101110110000111111011111011;
		correct = 32'b11011111111110011111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110011111101011001000101111;
		b = 32'b11011000110110110100001100101100;
		correct = 32'b11011110111111111111001100101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000100000111111000011101111;
		b = 32'b00011111001010011101111111000111;
		correct = 32'b10111111101010111111111111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011011101010101110110111010;
		b = 32'b01000000111001100101011101110101;
		correct = 32'b01001011111101110101111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110110010010011111000000100100;
		b = 32'b10001010110110011010100111001111;
		correct = 32'b11111110110110011111100111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000110110110011000000011001;
		b = 32'b11111111010111011001001010100111;
		correct = 32'b11111111110111111011001010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000100110110011110001101001;
		b = 32'b10010000011001110111000110110101;
		correct = 32'b11110000111111110111110111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111001101000010001011001101;
		b = 32'b11010101100111000100101111011101;
		correct = 32'b11111111101111000110101111011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001001010011110110001011111;
		b = 32'b10110000101110101000101000110111;
		correct = 32'b11110001101110111110111001111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100010100010001010101010001;
		b = 32'b10111100011101000110010000010011;
		correct = 32'b11111100011101010111010101010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110101000111110011000000010;
		b = 32'b00000100101011001100011000100001;
		correct = 32'b00110110101011111110011000100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000010100001001111111000000;
		b = 32'b10110000101110001110111011100011;
		correct = 32'b11110000111110001111111111100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010001000001001010010000001;
		b = 32'b01011101011101001001100110011110;
		correct = 32'b01111111011101001001110110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101111010111001101100100101;
		b = 32'b01110000111000000000010011111001;
		correct = 32'b01110101111010111001111111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100001010101000011000101100;
		b = 32'b00100001011000011111001010111011;
		correct = 32'b10100101011010111111011010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110101000001010111111001110;
		b = 32'b00100011011111100010010100100011;
		correct = 32'b01110111111111101010111111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000010011001001011011000110;
		b = 32'b01010100001101100110111001101010;
		correct = 32'b11010100011111101111111011101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010000100001110110110101000;
		b = 32'b00011100001100000100110100100100;
		correct = 32'b00111110001100001110110110101100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100001111111011111010111011;
		b = 32'b10111111010011011011101110101011;
		correct = 32'b11111111011111111011111110111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110011111011101000010100100;
		b = 32'b00000110101011101000010110110011;
		correct = 32'b00101110111111111101010110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110111111000011010101000001;
		b = 32'b11101100100110101011010100100110;
		correct = 32'b11101110111111101011010101100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100101100000010000111100111;
		b = 32'b11100011110110101110000010001001;
		correct = 32'b11100111111110101110000111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110000011111111001110001111;
		b = 32'b11000110011110110000101010111000;
		correct = 32'b11001110011111111111101110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000010000110011001100111001;
		b = 32'b01101111110111000101000100111100;
		correct = 32'b11101111110111110111001100111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101111001010000011100001011;
		b = 32'b01000100011010111010011110010100;
		correct = 32'b01010101111011111010011110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010110001101101101011111000;
		b = 32'b11101001100100100101011100011011;
		correct = 32'b11111011110101101101111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111100101010000011101001101;
		b = 32'b11000001101110101100011010010001;
		correct = 32'b11011111101111111100011111011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110101100111000010100100001;
		b = 32'b00010101100010100001110001111110;
		correct = 32'b00010111101110111001110101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010100111011100100110100100;
		b = 32'b01110010000110010001110101011000;
		correct = 32'b01110010100111011101110111111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000111000110011100001111111;
		b = 32'b11101100110110110111010111011111;
		correct = 32'b11111100111110110111110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011001000101100100010111100;
		b = 32'b01001000111011010111111010010100;
		correct = 32'b01011011111011111111111010111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111010100010010101110011111;
		b = 32'b00001101100000000010000011011001;
		correct = 32'b10111111110100010010101111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111101001011010100110011110;
		b = 32'b10100111001001101100011001111101;
		correct = 32'b10101111101001111110111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010100000010110001101000011;
		b = 32'b10010010010101011100011010111000;
		correct = 32'b11010010110101011110011111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110100001001000001011101011000;
		b = 32'b00011011101001010101110001111110;
		correct = 32'b10111111101001010101111101111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011111000100110111001111101;
		b = 32'b10111010100101110001111100000000;
		correct = 32'b10111011111101110111111101111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101110110011100100111100111;
		b = 32'b11111000111110100100110100111110;
		correct = 32'b11111101111110111100110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001011110001111110101010110;
		b = 32'b11001111111110010011111011000001;
		correct = 32'b11101111111110011111111111010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110001110110111010011001010;
		b = 32'b10100011101000101101100001100011;
		correct = 32'b11100111101110111111110011101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011110010010111000001110011;
		b = 32'b11101010001000001111001000110111;
		correct = 32'b11111011111010011111001001110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001101000100110110010010101;
		b = 32'b01011111111000111000011011011000;
		correct = 32'b01011111111000111110111011011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001101111001010100110101010;
		b = 32'b00000011111110011010010111010101;
		correct = 32'b11101011111111011010110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000011110110000000001101110;
		b = 32'b00111110010001010001110000011000;
		correct = 32'b10111110011111110001110001111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110010011101101010000010110;
		b = 32'b01000001110111101101100001001101;
		correct = 32'b01000111110111101101110001011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101100111101010001101100100;
		b = 32'b11010011110101101011100010000100;
		correct = 32'b11011111110111101011101111100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100010100100011111100100000;
		b = 32'b10010011000101111010110000100100;
		correct = 32'b10010111010101111011111100100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001100000111110101110010100;
		b = 32'b01101001010101011110001000111001;
		correct = 32'b11111001110101111110101110111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100100111000011110001011000;
		b = 32'b11000110100000011011100101110000;
		correct = 32'b11011110100111011011110101111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000001001000111100101110110;
		b = 32'b10000100001000100000011010100000;
		correct = 32'b11000100001001100111111111110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010111101111101010001111001;
		b = 32'b10100101011100111001010010101001;
		correct = 32'b10100111111101111101010011111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101011001001011010111100011;
		b = 32'b11110000011100000011111110110110;
		correct = 32'b11110101011101001011111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001101100001001011100100000;
		b = 32'b10001000011100110010100011011011;
		correct = 32'b10001001111100111011111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010011011111100110100100000;
		b = 32'b10111101111101101100011110011100;
		correct = 32'b11111111111111111100111110111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100101010011001100000101011;
		b = 32'b01101101011100100110110000101011;
		correct = 32'b11111101111110111111110000101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000101111000000010001101111;
		b = 32'b10110100101010110001110111000111;
		correct = 32'b11110100101111110001110111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011010110101011101001100100;
		b = 32'b10000001000010001011111111000011;
		correct = 32'b10101011010110101011111111100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110001101011000110000101101;
		b = 32'b11100001110110110101000100110001;
		correct = 32'b11110111111111111101110100111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010001100000000111010110100;
		b = 32'b11011110110000000110101110101110;
		correct = 32'b11011110111100000110111110111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110001111101100011100010011;
		b = 32'b11010110000001000101101110001100;
		correct = 32'b11110110001111101101111110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011010000011011001110110101;
		b = 32'b00100101100010110101011001001000;
		correct = 32'b11100111110010111111011111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101100000010000000001011110001;
		b = 32'b01111111010000100110100111100100;
		correct = 32'b01111111010010100110101111110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111000010000110100011101101000;
		b = 32'b10110001010001010100100011100000;
		correct = 32'b11111001010001110100111111101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100101110001110011000000011111;
		b = 32'b00010001010011111010101100010101;
		correct = 32'b01110101110011111011101100011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111101001011001000110101101;
		b = 32'b01101001001100111011010101100111;
		correct = 32'b01101111101101111011010111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011010000100011110101101000;
		b = 32'b10100011110110001010101000110101;
		correct = 32'b10110011110110101011111101111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110010101110101111101110010;
		b = 32'b11101010110110110000111110101001;
		correct = 32'b11111110110111110101111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110101001111100010101011001;
		b = 32'b11100100100111011101010000011101;
		correct = 32'b11110110101111111101010101011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100110010111111101110110101;
		b = 32'b10000110111111110110111010110010;
		correct = 32'b10010110111111111111111110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001110101100011110000001111;
		b = 32'b00000010100110101001011111000100;
		correct = 32'b10100011110111101011111111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100000111110001100000111110;
		b = 32'b00010011000011010010100011111001;
		correct = 32'b11010111000111110011100011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001101110101000100010001101;
		b = 32'b11110011110110100010100000110100;
		correct = 32'b11110011111110101010100010111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001000101010110101101010000;
		b = 32'b00111111010000111110001100100001;
		correct = 32'b01111111010101111110101101110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101100011100111000001101111;
		b = 32'b00100101010010101101011111111001;
		correct = 32'b11100101110011101111011111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110010101000001011000011010;
		b = 32'b01011110101010010101001110110101;
		correct = 32'b01011110111111010101011110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001010011011001100111100101;
		b = 32'b11110000100100101011001101010111;
		correct = 32'b11110001110111111011101111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000001001110000001000111011;
		b = 32'b00111101111011111111010100111110;
		correct = 32'b01111101111011111111011100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011011010010110000111101110;
		b = 32'b01000100010110010010100001100000;
		correct = 32'b01000111011110010110100111101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010110110110010100010100100;
		b = 32'b10001100011000011101000110010110;
		correct = 32'b10001110111110111111100110110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001111101110101001011010000;
		b = 32'b10000110110110010011011110100010;
		correct = 32'b11000111111111110111011111110010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011011110001101010001010011;
		b = 32'b11111111000111011101111000000011;
		correct = 32'b11111111011111011101111001010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011110000101111100111101001;
		b = 32'b00011100011010000010100001001110;
		correct = 32'b01111111111010101111100111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010110000000101110001100101111;
		b = 32'b01000010010111011110110111110000;
		correct = 32'b11010110010111111110111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101011111110001110011001110;
		b = 32'b10000011010011011010011001001000;
		correct = 32'b10110111011111111011111011001110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101010111010000111000101101;
		b = 32'b00010001111101010101110001101000;
		correct = 32'b01011101111111010101111001101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011010100000110000000100100;
		b = 32'b11101110011011001111011010001001;
		correct = 32'b11111111011111001111011010101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100011111011001110101100000110;
		b = 32'b01100001001000101110111111111111;
		correct = 32'b01100011111011101110111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011110000011111001010111000;
		b = 32'b10001011010000011001100101001001;
		correct = 32'b11111011110000011111101111111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010101001001000111110000110;
		b = 32'b11001101001001100011101101010101;
		correct = 32'b11011111101001101011111111010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000001000000100010111110100;
		b = 32'b10001100011101011000111001101111;
		correct = 32'b10011100011101011100111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001101110110101100001110001;
		b = 32'b01010100110011111101010101011101;
		correct = 32'b11111101111111111101110101111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010000010101000001011000111;
		b = 32'b10000100111011010111101011000000;
		correct = 32'b11011110111011111111101011000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000101000110110100000001010;
		b = 32'b10101000011000011010101101110110;
		correct = 32'b11111000111000111110101101111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010010010101010111010110100;
		b = 32'b00111001111100110110001011011111;
		correct = 32'b00111011111110111110111011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001010000001100111111010011;
		b = 32'b10110101111010110011010001001110;
		correct = 32'b11110101111010111111111111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100101001110010010111000110;
		b = 32'b00000101000110011011100101100101;
		correct = 32'b10100101101111111011110111100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110001110111111101010001110;
		b = 32'b01100101111010010000101000100111;
		correct = 32'b01111111111110111111101010101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010000110100000011001101001;
		b = 32'b00101111111111111010100000011100;
		correct = 32'b10101111111111111010111001111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001010000010111111111101010;
		b = 32'b00101000001000100011100000000001;
		correct = 32'b11111001011000110111111111101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110101100111011011011000000;
		b = 32'b10001111000110111011110101100111;
		correct = 32'b10111111101110111011111111100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000000101011000100010100001;
		b = 32'b10011101100011100101000101000110;
		correct = 32'b11011101100111111101100111100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011011100000110001001110000;
		b = 32'b00010111101111011101001010110011;
		correct = 32'b01010111111111011111001011110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000110110110010101010011100;
		b = 32'b01010111100011101000101111011110;
		correct = 32'b01110111110111111010101111011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110111100000100110000011111;
		b = 32'b11000010110010101000110100100001;
		correct = 32'b11011110111110101100110100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011011101000000000001110100;
		b = 32'b00111011011110101010110010010101;
		correct = 32'b10111011011111101010110011110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111101110100110111001111010;
		b = 32'b00000000101100111010101010011100;
		correct = 32'b11001111101110111110111011111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100000100010100000000011010;
		b = 32'b00010101101100100001010010101010;
		correct = 32'b00011101101100110101010010111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001101101101110111011011001011;
		b = 32'b01110011001100101110101001001101;
		correct = 32'b01111111101101111111111011001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101010010111110000101001111;
		b = 32'b11100011110010001101000111110110;
		correct = 32'b11101111110010111111000111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100011100001001111110100110;
		b = 32'b01100010110011001111001010001111;
		correct = 32'b01110110111111001111111110101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000110011001011111000011011;
		b = 32'b11101111010011110100011100010111;
		correct = 32'b11111111110011111111111100011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000110110000010011110100101;
		b = 32'b10010110101001000111111111111011;
		correct = 32'b11010110111111000111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101000000011111110001110100;
		b = 32'b10001111111000111100001110101110;
		correct = 32'b11111111111000111111111111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100110010101010001111111001;
		b = 32'b11111101111111000110101110101000;
		correct = 32'b11111101111111101110101111111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111010100111110010110101010;
		b = 32'b00000110111011011010010101101110;
		correct = 32'b11000111111111111110010111101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011000011101000101110011100;
		b = 32'b11010110000000110100001110111010;
		correct = 32'b11010111000011111100101110111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011010010010111110100010011;
		b = 32'b01101101110110000110000101100110;
		correct = 32'b01111111110110010111110101110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010001100000111001001101101;
		b = 32'b10110001100101000101011110000110;
		correct = 32'b10110011101101000111011111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001010110000011001010011011;
		b = 32'b10010000100011000000011101001011;
		correct = 32'b10011001110111000011011111011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110010001110101000000000010;
		b = 32'b01110010001101101101111011011111;
		correct = 32'b01110110011101111101111011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101111011111000011101000001;
		b = 32'b01100001001110110010111110000010;
		correct = 32'b11110101111111111010111111000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100100011100000101000011101;
		b = 32'b10011110100100110001000101000011;
		correct = 32'b11011110100111110001101101011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100011111110010011011111000;
		b = 32'b10001011010101101100110110010001;
		correct = 32'b10001111011111111110111111111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110000111111011011110101111;
		b = 32'b01111111110010001001111101010010;
		correct = 32'b11111111110111111011111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101001101001100101011000100;
		b = 32'b00000101111101110100010111110010;
		correct = 32'b11001101111101111100111111110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101111001001001110010001000;
		b = 32'b10111010000101000001011110101000;
		correct = 32'b10111111111101001001111110101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111111110010010010101000111;
		b = 32'b11001010101001110110000101001100;
		correct = 32'b11001111111111110110010101001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010111011001101011000111011;
		b = 32'b00011000111101101111100001011110;
		correct = 32'b00111010111111101111111001111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100110010100001001010010111;
		b = 32'b11110110100000101111100011010000;
		correct = 32'b11110110110010101111101011010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001011110011111001000000111;
		b = 32'b10001000010000111101111011011110;
		correct = 32'b10001001011110111111111011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011101010001110011100111101;
		b = 32'b00000000101001101110000010010111;
		correct = 32'b11001011101011101110011110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000001010101010110100110001;
		b = 32'b11111100101111011101111101100101;
		correct = 32'b11111100101111111111111101110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011110001100110010110001011;
		b = 32'b11000010100110000100111001110011;
		correct = 32'b11010011110111100110111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110101000110101111100100010;
		b = 32'b10000010101111100100001000010011;
		correct = 32'b10110110101111110101111100110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011111101111111111101000011;
		b = 32'b11001110110001010001101101000100;
		correct = 32'b11011111111101111111111101000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000010110001110011000000011;
		b = 32'b01010110010011011110011110111101;
		correct = 32'b01011110010111011110011110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101101100101110111101001001;
		b = 32'b00000000110011100101011000001001;
		correct = 32'b00100101111111101111111101001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101000110100011011101100110;
		b = 32'b11001011110011011001010100101001;
		correct = 32'b11101111110111111011011101101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001001111010011001100100110;
		b = 32'b11011001010000110000110010110101;
		correct = 32'b11011001011111110011111110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001101111010111101101110101;
		b = 32'b01000101101010001001001001000010;
		correct = 32'b11101101101111011111101101110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100001111001100111011110111;
		b = 32'b00100010100101010101101010101010;
		correct = 32'b00100110101111011101111011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011110110101111111101100011;
		b = 32'b10011001001100100111100000100001;
		correct = 32'b10011011111110101111111101100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011101010001111100110101001;
		b = 32'b00111110100110000010100001111010;
		correct = 32'b01111111101110001111100111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111110000110111011110011011;
		b = 32'b10010110011010000110110000001000;
		correct = 32'b10110111111010110111111110011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100010000001101011001001111;
		b = 32'b10010110110111010111011011100100;
		correct = 32'b10011110110111011111011011101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101000011101101101100011101;
		b = 32'b01010000001111101010101001011100;
		correct = 32'b11011101001111101111101101011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101001000100010110010111011;
		b = 32'b01101100011010001010111101011011;
		correct = 32'b11101101011010101010111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011000100010100001011100100;
		b = 32'b10011011001110101000111100000010;
		correct = 32'b11111011001110111100111111100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001101101000110001001111011;
		b = 32'b00010010010001100100111011000110;
		correct = 32'b01111011111101100110111011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000110111011111110011000100;
		b = 32'b01011110011111001111100111000100;
		correct = 32'b01111110111111011111110111000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010011101110111011110000000;
		b = 32'b00000010100101100100100011010001;
		correct = 32'b10100010111101110111111111010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110111101000011010100110111;
		b = 32'b01100111100000011011000011000101;
		correct = 32'b01101111111101011011010111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000111011011101101000100101;
		b = 32'b00111111011100000010010010001000;
		correct = 32'b11111111111111011111111010101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010101011100100010110011001111;
		b = 32'b11011000101100111001100100010101;
		correct = 32'b11011101111100111011110111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010111011110001010100000110;
		b = 32'b10001110111110011011001000110110;
		correct = 32'b11101110111111111011011100110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011010101100001111101001010;
		b = 32'b00110000101001110011011100111001;
		correct = 32'b11110011111101110011111101111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110011000110100100101101010;
		b = 32'b00001011101111111011110000110101;
		correct = 32'b11101111111111111111110101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011001000001100100010111111;
		b = 32'b00111000101001011111010001101000;
		correct = 32'b01111011101001011111110011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101001011001001011100100101;
		b = 32'b10010000011010000100110110101000;
		correct = 32'b11110101011011001101111110101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110110011000110001100001000;
		b = 32'b11010100011000000100011010011100;
		correct = 32'b11010110111011000110011110011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011110111001010001011100111;
		b = 32'b01110111001101001001101000010100;
		correct = 32'b01111111111111001011101011110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010011010111001000001010011;
		b = 32'b00000011000100010110001001101001;
		correct = 32'b10111011011110111111001001111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011001111001000100001111000;
		b = 32'b00000010100011011000000010011010;
		correct = 32'b01111011101111011000100011111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000000100111011011100000110;
		b = 32'b01111011010101011111011100111001;
		correct = 32'b01111011010101111111011100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100100111101110010111100000;
		b = 32'b11000111100000011001111111110101;
		correct = 32'b11100111100111111111111111110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011100100010010010101100101;
		b = 32'b00001101111010000101011000001111;
		correct = 32'b01101111111110010111011101101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101010111111010010001001000;
		b = 32'b01111000101111011001001111000000;
		correct = 32'b11111101111111111011011111001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111011110111001011000011100;
		b = 32'b11010000000010011110101111010011;
		correct = 32'b11011111011110111111111111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001101000010110011110011000;
		b = 32'b10111101011011111010001011111000;
		correct = 32'b10111101111011111110011111111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011111101010101011001010000;
		b = 32'b01101111011111010110001000100000;
		correct = 32'b01111111111111010111011001110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000000011101110010010000010;
		b = 32'b01100001011101110100111010010011;
		correct = 32'b01101001011111111110111010010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110110100011110111001110110;
		b = 32'b10000101110100110100010001000101;
		correct = 32'b11010111110100111110111001110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100100000010111100001000001000;
		b = 32'b01000111001010110001111111101010;
		correct = 32'b01100111001010111101111111101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011011010001100010101011110;
		b = 32'b11000010011100010001100000000110;
		correct = 32'b11011011011110011101110101011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101001110110010010001010101;
		b = 32'b01100111110011011101100001001011;
		correct = 32'b01111111111111111111110001011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011111001101110111000100000;
		b = 32'b01001110101001101001001000010000;
		correct = 32'b11001111111001101111111000110000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110010110010101111011000110;
		b = 32'b10001001110101111001010110100001;
		correct = 32'b11101111110111111101111111100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100010110111101000011101100;
		b = 32'b11011001110010111000011100101111;
		correct = 32'b11011101110110111101011111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000101000101010100010011001;
		b = 32'b10100111001100110100001010110011;
		correct = 32'b10110111101100111110101010111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110010010001010001010110001;
		b = 32'b00100001100101101000000101101111;
		correct = 32'b10101111110111101010001111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010000110111001111010001111;
		b = 32'b10110101000100101110001110001010;
		correct = 32'b11110111000110111111111110001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100010110100101001100010000;
		b = 32'b00111101000000100001101110000010;
		correct = 32'b10111101010110100101101110010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100111000110111010110100100011;
		b = 32'b00101011011100010001001010101101;
		correct = 32'b00101111011110111011111110101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010111111101101111110001001;
		b = 32'b01001000110100100010101111001111;
		correct = 32'b01001010111111101111111111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010001100011000011001100110;
		b = 32'b00101100110000010011011110100000;
		correct = 32'b01111110111100011011011111100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000001101000110010111100101;
		b = 32'b10111011111011101101000111001010;
		correct = 32'b11111011111111101111010111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001101011111100011001010110;
		b = 32'b11001110101000111001110100110110;
		correct = 32'b11111111101011111101111101110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110111000001001110000011001000;
		b = 32'b11000111111010000111011101111100;
		correct = 32'b11110111111011001111011111111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000111101100001000100001010;
		b = 32'b00100011100110101110101111110110;
		correct = 32'b00111011111111101111101111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111110010110101001101001001;
		b = 32'b00000101000000011110110011011111;
		correct = 32'b01001111110010111111111111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001011000000101101101010011;
		b = 32'b00010001110101101000110010101010;
		correct = 32'b00110001111101101101111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101011101111010101111111100;
		b = 32'b11001000011010101011101010100011;
		correct = 32'b11111101011111111011101111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101000011101110110110100010;
		b = 32'b00101000111101001011110011010011;
		correct = 32'b00111101111111101111110111110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010110000011011011001100101;
		b = 32'b11000000010010010001100001011001;
		correct = 32'b11000010110010011011111001111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101110010100010101100111111;
		b = 32'b11001010100010000101011010000011;
		correct = 32'b11011111110010100111111110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010000101110000010111111000;
		b = 32'b10010011011010100101011010010100;
		correct = 32'b10010011011111110101011111111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110000001110100011110001111;
		b = 32'b10011000010100111001011010001010;
		correct = 32'b11111110010101111101011110001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011101000000100000111011110;
		b = 32'b11101010111100111010001101010001;
		correct = 32'b11101011111100111110001111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101001101111011000011101001;
		b = 32'b01111100001000110101100100011000;
		correct = 32'b01111101001101111111100111111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001100111000011000101001000;
		b = 32'b10010011110111010000101011000100;
		correct = 32'b10010011110111010011101111001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001011110100010111011100111;
		b = 32'b10100110110011010100110111010000;
		correct = 32'b11100111111111110110111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111000101100001100101100111001;
		b = 32'b00100010010101001011111111000110;
		correct = 32'b11111010111101001111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010100010000100000011111100;
		b = 32'b10111101111100110111010010100010;
		correct = 32'b10111111111110110111010011111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110010000011011101001011000;
		b = 32'b00011110111001110111111100000000;
		correct = 32'b00011110111001111111111101011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100011011010110110111010000;
		b = 32'b11101011110111100010100001101011;
		correct = 32'b11101111111111110110110111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001011010101110111001001010;
		b = 32'b10001111011000000101000000110001;
		correct = 32'b10001111011010101111111001111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111010000110011110111101001;
		b = 32'b00110111001101110110100011000001;
		correct = 32'b00110111011101110111110111101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111101011001011001010101110;
		b = 32'b00010010101111110011101101101001;
		correct = 32'b01111111101111111011101111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010111011111110011110001111;
		b = 32'b00100101011101011010110000010011;
		correct = 32'b10111111111111111110111110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000001110010000001001100011111;
		b = 32'b11110001100011001001101011011100;
		correct = 32'b11110001110011001001101111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111110001000110100101010000;
		b = 32'b10011101110101100110101011111000;
		correct = 32'b10111111110101100110101111111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010101001111001011000011110;
		b = 32'b01010101001000100011101110011010;
		correct = 32'b01110111101001111011111110011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100110100010111001110111101;
		b = 32'b11101010111111001000000110011011;
		correct = 32'b11101110111111011111001110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111011101110011110010011001;
		b = 32'b00010110001001000001010111100101;
		correct = 32'b01110111011101110011110111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000110101111010011001000100;
		b = 32'b00001111100110111111001110010010;
		correct = 32'b00101111110111111111011111010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110100100000001101001110110;
		b = 32'b00100110000110110000101111010111;
		correct = 32'b10110110100110110001101111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111111000110001011100000111;
		b = 32'b01010100110010000110010101100001;
		correct = 32'b01111111111010110111011101100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010001001101100101110010010;
		b = 32'b01110101010011101111101001110111;
		correct = 32'b01111111011011101111101111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111011011001000011010101011;
		b = 32'b00000010000111011010001100100010;
		correct = 32'b10110111011111011010011110101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000100000100110011001010101010;
		b = 32'b11011111001110000001100111011011;
		correct = 32'b11011111001110110011101111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100001101111111011001100000010;
		b = 32'b00000011111101101111001110010000;
		correct = 32'b00100011111111111111001110010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111010011001101011110100101;
		b = 32'b10111010101110110101101001110000;
		correct = 32'b10111111111111111101111111110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000100100111010001101000111;
		b = 32'b00101101110001010101110101100111;
		correct = 32'b01101101110101111111111101100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110101110101100100010001110;
		b = 32'b10010111010011111101101111111111;
		correct = 32'b10111111111111111101101111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110010100101010100111101011;
		b = 32'b11100011111111000000001101100111;
		correct = 32'b11100111111111101010101111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101111100000000101111010001;
		b = 32'b00011100010110001011111001100011;
		correct = 32'b11111101111110001011111111110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110011000100011000001011000;
		b = 32'b11111011111100100110011000101100;
		correct = 32'b11111111111100100111011001111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101011100010111100111011111;
		b = 32'b00110111000101100100000010101001;
		correct = 32'b00110111011101110111100111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111011110101001010000011011;
		b = 32'b00111101101001101011010111000001;
		correct = 32'b01111111111111101011010111011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101000101000101010000100100;
		b = 32'b11101001010111101111110101111100;
		correct = 32'b11111101010111101111110101111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010001100111100001100101100;
		b = 32'b00101000010011001110011110111100;
		correct = 32'b10111010011111111110011110111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110110110110011010010100000;
		b = 32'b11001000110111100011100111111111;
		correct = 32'b11101110110111110011110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000011000011010111011001001;
		b = 32'b11000110110101001111110000111011;
		correct = 32'b11000110111101011111111011111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001111000010001101110000010;
		b = 32'b10101001111000000100000110011010;
		correct = 32'b11101001111000010101101110011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100001011000100110101000010;
		b = 32'b10100010110001101110011011010110;
		correct = 32'b10101110111011101110111111010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010000000010001001011100101;
		b = 32'b11111111000000001011111100110011;
		correct = 32'b11111111000000011011111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011100111111000110001000110;
		b = 32'b01101010011010001010000000101001;
		correct = 32'b11101011111111111010110001101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010001110001110010000111010;
		b = 32'b11000111010000111110101111001101;
		correct = 32'b11011111011110111110111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101111101000110010001100111;
		b = 32'b00000111110110111001100100110101;
		correct = 32'b01101111111111111111110101110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110010000101000000110100100;
		b = 32'b00011001000101000000011000011111;
		correct = 32'b00111111010101101000011110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101111011101011101000100110;
		b = 32'b01011110101100000100101000010011;
		correct = 32'b11011111111111101111101000110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100101111100100011101000100;
		b = 32'b11101101001111110100011010101101;
		correct = 32'b11101101101111110100011111101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010101111110000111101110000;
		b = 32'b01001011110011100111010000100010;
		correct = 32'b01101011111111110111111101110010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000100000011001010000001100010;
		b = 32'b01110000101100101000111010001000;
		correct = 32'b11110100101111101010111011101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001110100011011010001100001;
		b = 32'b11011000010001011001101001110001;
		correct = 32'b11011001110101011011111001110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101101000100101001110111011;
		b = 32'b01110011000010010110000001001011;
		correct = 32'b11111111101010110111001111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000010010010100000101011011;
		b = 32'b11111011010010101110111110110011;
		correct = 32'b11111011010010111110111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100001010011011101101001101;
		b = 32'b01000111011110110110110010111011;
		correct = 32'b11010111011110111111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101011100101100100110110010;
		b = 32'b10101110110101000001011110010011;
		correct = 32'b11111111111101101101111110110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011111011001111100000011000;
		b = 32'b11010000101010110010101010101000;
		correct = 32'b11110011111011111111101010111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011010011000110001001001000;
		b = 32'b01010111110010101110100010001000;
		correct = 32'b01110111110011101110101011001000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110010011000100001011111111;
		b = 32'b01011001001100010001101010101000;
		correct = 32'b11111111011111010101101011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101101001010001001101000001;
		b = 32'b00010100110001101100110001100111;
		correct = 32'b01111101111001111101111101100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101001011111100111011110000;
		b = 32'b01011001000110001100110111011000;
		correct = 32'b01111101001111111100111111111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100001000010000000110111000110;
		b = 32'b11101001001010111010000110010011;
		correct = 32'b11101001001010111010110111010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011110010101110110101001011;
		b = 32'b00101100101000110111100001000101;
		correct = 32'b11101111111010111111110101001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101000100000000010100000011;
		b = 32'b10010101000010000100000110110101;
		correct = 32'b11111101000110000100010110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011010101110101100111110010;
		b = 32'b00001001010100101010110110100111;
		correct = 32'b00001011010101111111110111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010010101111111111111010011;
		b = 32'b10000100110110000010010001010011;
		correct = 32'b10010110110111111111111111010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001010111000010100100110111;
		b = 32'b01110101101001011010011101000001;
		correct = 32'b11110101111111011010111101110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010110010100110100000000110;
		b = 32'b01111011010100110001110001111001;
		correct = 32'b01111011110110110111110001111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010110111000110111010111110;
		b = 32'b01001111100100010100110101101110;
		correct = 32'b11101111110111010110111111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101011001101010100011000100000;
		b = 32'b01101011011001110010001111010110;
		correct = 32'b11101011011101110110011111110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010011001101101101101100100100;
		b = 32'b11101110101000000010000101100001;
		correct = 32'b11111111101101101111101101100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110111011101101000011011110;
		b = 32'b00010101100010000111011000100011;
		correct = 32'b00110111111011101111011011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000110001101001001101011110;
		b = 32'b01101110110110100011101101010010;
		correct = 32'b01111110110111101011101101011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101111010000000010000000111011;
		b = 32'b00110000010101110010111011111010;
		correct = 32'b11111111010101110010111011111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101110010000010111011100110;
		b = 32'b00010010011001001100011110110011;
		correct = 32'b11111111111011001110111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111000101101001101100101000;
		b = 32'b00101110110000000001010000011000;
		correct = 32'b11101111110101101001111100111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010100110011110011101100101;
		b = 32'b00100010000000111111010100011100;
		correct = 32'b00111010100110111111011101111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000110011011110101010100011;
		b = 32'b10110000000101111010100000000110;
		correct = 32'b11111000110111111110101010100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111011000110111010100000111;
		b = 32'b01101111000110110111001010110111;
		correct = 32'b11101111011110110111011110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000100001010101110010010111100;
		b = 32'b00110110111011110101110011001000;
		correct = 32'b10110110111011111111110011111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011010111110010110011000100;
		b = 32'b01011010001010001101000011010001;
		correct = 32'b11011011011111111111110011010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110010111110001100101011100;
		b = 32'b01001110100010101011011100000011;
		correct = 32'b01111110110111111011111101011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111101000111001001011110000;
		b = 32'b11011010001100001000100000111110;
		correct = 32'b11011111101100111001101011111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100000010001010001010010000;
		b = 32'b11010010101100010111110111010110;
		correct = 32'b11011110101110011111111111010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010100100100111010011100001;
		b = 32'b01100111110110110010001111101011;
		correct = 32'b01111111110110110111011111101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100001011101100001011010001;
		b = 32'b11100000101001101111101011000110;
		correct = 32'b11110100101011101111101011010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000100000110011101011101011;
		b = 32'b11000011010010111011101101111010;
		correct = 32'b11000011110010111011101111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011110111101001111010011100;
		b = 32'b01100010100111111011001011100100;
		correct = 32'b11111011110111111011111011111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001010011010100110101111000;
		b = 32'b01011010010110101100011110110001;
		correct = 32'b11111011010111111100111111111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000111101001101011010111000;
		b = 32'b11100111101111110001010101001011;
		correct = 32'b11101111111111111101011111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011111001110011011010000000;
		b = 32'b10011011011110100111011101100010;
		correct = 32'b11011011111111110111011111100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110110101100011100000101001;
		b = 32'b00101010111000100010111000110100;
		correct = 32'b00111110111101100011111000111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001000010011111000101010011;
		b = 32'b10100101100111011011110000110000;
		correct = 32'b10111101100111011111110101110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101111000111110111110010110;
		b = 32'b01111001100101100001101101111011;
		correct = 32'b01111101111101111111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000100110100100111110000011;
		b = 32'b11110101100001111010111010001101;
		correct = 32'b11111101100111111110111110001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010110001110001001010100010;
		b = 32'b00010110100111010111101111000011;
		correct = 32'b01010110110111110111101111100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110101011010110100001001011000;
		b = 32'b11000111001011100011111000111111;
		correct = 32'b11110111011011110111111001111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001100111111101010100101110010;
		b = 32'b00111010110000101110001011000011;
		correct = 32'b10111110111111101110101111110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101011110010101101110001110100;
		b = 32'b01001110000101100101000010101001;
		correct = 32'b11101111110111101101110011111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111101000111101111000110110;
		b = 32'b10001101101011100011100111110001;
		correct = 32'b11111111101011111111111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011011110100011010110000111;
		b = 32'b10001011110010111100101100010100;
		correct = 32'b10011011111110111111111110010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110010100000110001110011100;
		b = 32'b10100011000010100000110000011111;
		correct = 32'b10101111010110100110111110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011001010011001111110100011;
		b = 32'b10011111100001011111100001010011;
		correct = 32'b10111111101011011111111111110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110111011101011010001001010;
		b = 32'b10110011010101010111110110010100;
		correct = 32'b11111111111111111111110111011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110110010011001000100010011100;
		b = 32'b11110001010001110001010101001000;
		correct = 32'b11110111010011111001110111011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101101011011111111000011101;
		b = 32'b11111101000001100011111111010101;
		correct = 32'b11111101101011111111111111011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110000101000000110110001110;
		b = 32'b11010111101011100001011000101111;
		correct = 32'b11110111101111100001111110101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000100010011101111101110100;
		b = 32'b01110011101011000101011100011100;
		correct = 32'b01111011101011011101111101111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011111100101001111110001001;
		b = 32'b00111111001101100110000000010011;
		correct = 32'b10111111111101101111111110011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000111101000101010111000001;
		b = 32'b01100011010001000011001110110010;
		correct = 32'b01110011111101000111011111110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111001111100000101011110000;
		b = 32'b01010011001001101100100000100101;
		correct = 32'b11010111001111101100101011110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011100111000000101000100110;
		b = 32'b00000001001101011110111011000111;
		correct = 32'b10000011101111011110111011100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010000101111110011100010010;
		b = 32'b11001010110010111110100011100111;
		correct = 32'b11111010110111111110111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100101101011010010110110111;
		b = 32'b01010101001101110011011111111001;
		correct = 32'b11010101101101111011011111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000000000010101110100101111;
		b = 32'b10001000111111100010101011100110;
		correct = 32'b11011000111111110111111111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011010110110011010101011010;
		b = 32'b11000100011100110111100000111011;
		correct = 32'b11010111011110110111110101111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001111101100001011101110101;
		b = 32'b00010011100100011010001110110100;
		correct = 32'b10110011111101111011011111110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000000100010111101001010001;
		b = 32'b00101001001100111000001001101111;
		correct = 32'b11101001001100111111101001111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000110101000111010001100010;
		b = 32'b00111100001011011101110101110111;
		correct = 32'b10111100111111011111110101110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011101000100100110010101110;
		b = 32'b01111100011000100101000101110101;
		correct = 32'b01111111111000100101110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101000000100101101111110101;
		b = 32'b10001011110100010000000110010101;
		correct = 32'b10101111110100110101101111110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011111000110100100111011111;
		b = 32'b10010000101101011111101011010110;
		correct = 32'b10011011111101111111101111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111101111000110111010101101101;
		b = 32'b01100001111011100101011100011111;
		correct = 32'b01111101111011110111011101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111100011101100111111010010;
		b = 32'b01110000101101011110101111110111;
		correct = 32'b11111111101111111110111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111001000100001001111000100;
		b = 32'b11010110010011000011000111000110;
		correct = 32'b11011111011011100011001111000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100010010111101010000010110011;
		b = 32'b11001100011010011010101110100100;
		correct = 32'b11101110011111111010101110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111111110101011110111000001;
		b = 32'b01101100010011001011111011100011;
		correct = 32'b01111111111111101011111111100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010100100111110101001111110110;
		b = 32'b11011100000101110100011100001010;
		correct = 32'b11011100100111110101011111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101110010011011001010110001;
		b = 32'b01100111010010111010001011001101;
		correct = 32'b11111111110010111011001011111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010000111001111011111001110;
		b = 32'b01110100010100111000001100101100;
		correct = 32'b11111110010111111111011111101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000001101010101000010111010000;
		b = 32'b00010110011001001010001010011011;
		correct = 32'b00010111111011101010011111011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010100100110011111100001111;
		b = 32'b10011111100001011100110000010010;
		correct = 32'b10011111100101111111111100011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111110100100101010010000111;
		b = 32'b10001011110110011001110010010000;
		correct = 32'b10111111110110111101110010010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101101001101000000001101101;
		b = 32'b00100110000111101110011110011001;
		correct = 32'b10111111101111101110011111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111110001101110000000101100;
		b = 32'b10110100011100110001001010010111;
		correct = 32'b11110111111101111111001010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011000001000111111000000010;
		b = 32'b00101011001011001010111001111010;
		correct = 32'b11101011001011001111111001111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000110010110101100000010000;
		b = 32'b01001001110110100011011000011111;
		correct = 32'b01111001110110110111111000011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110010111011010010110011001;
		b = 32'b01100001001100111010111111000100;
		correct = 32'b11110111011111111010111111011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100010100111101011101000101;
		b = 32'b11111111111010111100000010001110;
		correct = 32'b11111111111110111101011111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101111001101100010011010000;
		b = 32'b01100001000100000010010000010101;
		correct = 32'b11100101111101101110010011010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100010000001010100101001100;
		b = 32'b10110111000100100101111101000101;
		correct = 32'b11110111010100101111111101001101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100011000110111011011000011;
		b = 32'b01010100111110100001100001001110;
		correct = 32'b01010100111110110111111011001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110010011011010100101011110;
		b = 32'b00010110101101111000010101010011;
		correct = 32'b00110110111111111010110101011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101010100010101001011100111;
		b = 32'b00100001100100111010101110110100;
		correct = 32'b11100101110100111111101111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111000101010110000101011000001;
		b = 32'b11010110000011000010111011010001;
		correct = 32'b11111110101011110010111011010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011111110100110100000011001;
		b = 32'b11101100100111010110110010010111;
		correct = 32'b11101111111111110110110010011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001010110001110000110011100;
		b = 32'b10001100101110101111011111101000;
		correct = 32'b11111101111110101111011111111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101001001111101111101011110;
		b = 32'b01011011110010000011101101111001;
		correct = 32'b01111111111011111111111101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101111100000101111000110110;
		b = 32'b01111110010001111110011111111110;
		correct = 32'b11111111111101111111111111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111011110010001000001000010;
		b = 32'b10010001101001011100000001111011;
		correct = 32'b11010111111111011101000001111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010000010100110101110010101000;
		b = 32'b11110000110010110110000001110111;
		correct = 32'b11110000110110110111110011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011101000001011010011011011;
		b = 32'b01100101011101101100110010110000;
		correct = 32'b01110111111101101111110011111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011110010100010110111100000;
		b = 32'b10001001010100010100111110110100;
		correct = 32'b11111011110110110110111111110100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000001110101110011010110101101;
		b = 32'b11010011111011010011010001101001;
		correct = 32'b11010011111111110011010111101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010110100100001000010010100;
		b = 32'b00010100011001100111110101010010;
		correct = 32'b00011110111101100111110111010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010001001000000111101111100;
		b = 32'b11110011111100111100011110010001;
		correct = 32'b11110011111101111100111111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101011100100001100101100110;
		b = 32'b11100010100011000111000111001111;
		correct = 32'b11110111111111100111100111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101010101001001010111110000;
		b = 32'b00100000001000011111100001010111;
		correct = 32'b01100101011101011111110111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101010010101000010111001010;
		b = 32'b10001010101111110010001111111100;
		correct = 32'b10011111111111111010011111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000000010110001011000010111;
		b = 32'b11101010101100110100000011101111;
		correct = 32'b11101010101110110101011011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100110100100110101010110111;
		b = 32'b00000100001110011001000011110001;
		correct = 32'b11111100111110111111101011110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010001101001110111101100111;
		b = 32'b00001111000011011101111010010000;
		correct = 32'b00101111001111011111111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110101010100101101010000101;
		b = 32'b10000100100111101100001000110011;
		correct = 32'b11101110101111101101101010110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100110101110011010101111001;
		b = 32'b01111111111011000011100100000010;
		correct = 32'b11111111111111110011110101111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111011100000011001001001001;
		b = 32'b01001100011101111011000100010010;
		correct = 32'b01111111011101111011001101011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110101110100111010100001101101;
		b = 32'b11110101011110010001101100111110;
		correct = 32'b11110101111110111011101101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010100110001010100100011001;
		b = 32'b01110001010100000000100101100010;
		correct = 32'b11110011110110001010100101111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111000101000011000011001100;
		b = 32'b00001001011111001100010101100111;
		correct = 32'b01001111011111001111010111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000010011011111001111101011;
		b = 32'b00101100000111011110110111000010;
		correct = 32'b10101100010111011111111111101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111111010101010100001100110;
		b = 32'b10011000100101110111011101010010;
		correct = 32'b11011111111111111111111101110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011111010110101010100101101;
		b = 32'b01001100101101010111001000010000;
		correct = 32'b11001111111111110111011100111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110000110000110111001011111;
		b = 32'b10110010101011011111011011011010;
		correct = 32'b10111110101111011111111011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101010110000101010110000010;
		b = 32'b00000111010111100110111101110110;
		correct = 32'b11010111010111100111111111110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000101110101011111100000011;
		b = 32'b11110111111001000010011100101011;
		correct = 32'b11110111111111101011111100101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000111011000100111010010011;
		b = 32'b11110100011110010110110001000011;
		correct = 32'b11110100111111010110111011010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110001110100111100010011110;
		b = 32'b10011111010101111001011111110101;
		correct = 32'b11111111011111111111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000101000110100100001000000001;
		b = 32'b01100100100110011111010100110100;
		correct = 32'b11100101100110111111011100110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110001101110101000011110101;
		b = 32'b00110011110001110000110110011000;
		correct = 32'b01111111111101110101110111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111010100111001011001100001;
		b = 32'b01100010010100111010101001101001;
		correct = 32'b11111111010100111011111001101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010010100000010000110101101;
		b = 32'b01100110101010011001000110111010;
		correct = 32'b01111110111110011011000110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010000011100111011111111000;
		b = 32'b11011100011111011011111100010111;
		correct = 32'b11111110011111111111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000000010110100110100111101010;
		b = 32'b10101011111111001010001111000001;
		correct = 32'b10101011111111101110101111101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001110101011111010011011100;
		b = 32'b11100011110001101001110100111110;
		correct = 32'b11110011110101111111110111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110101000011001001101100011001;
		b = 32'b00001010101111100100100011010011;
		correct = 32'b01111111101111101101101111011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111100100111011110111000101;
		b = 32'b10010111001101100100000100011011;
		correct = 32'b10011111101101111111110111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011111001100001000101111000010;
		b = 32'b00001111000100110101111011010011;
		correct = 32'b00011111001100111101111111010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011101011111010101100011101111;
		b = 32'b00110000111111101111100101010111;
		correct = 32'b01111101111111111111100111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110001111000000101011101111;
		b = 32'b01011101011100001100000100111100;
		correct = 32'b11111111011111001100101111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001110000011110111001101011;
		b = 32'b10001110100011110111000110010010;
		correct = 32'b11111111110011111111111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010010100101110110010011011001;
		b = 32'b10110100100001001001110001010011;
		correct = 32'b11110110100101111111110011011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111000101101110001010111000;
		b = 32'b11011100010000000011010101001010;
		correct = 32'b11011111010101101111011111111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110001000000111000110110011;
		b = 32'b10010011001111010000000110010110;
		correct = 32'b11111111001111010111000110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111011001000001010100111101;
		b = 32'b10111101111111100111110110000111;
		correct = 32'b11111111111111100111110110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110011010010000111001101111;
		b = 32'b01010000101001001011010101100001;
		correct = 32'b01110110111011011011111101101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111100101111111111011000111;
		b = 32'b00011001100010001001010100110000;
		correct = 32'b00011111100111111111111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110010000011001011000011010;
		b = 32'b00111100100111011000111011101100;
		correct = 32'b10111110110111011001111011111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001010110110110110111011111;
		b = 32'b11000100101000110010010100110011;
		correct = 32'b11001101111110110110110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011110000001000001101001101;
		b = 32'b10110110010001110010101010001011;
		correct = 32'b11111111110001111010101111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100001011010110001001010101;
		b = 32'b01010001100000011011111010111100;
		correct = 32'b01011101101011011111111011111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110101111101001011111101011;
		b = 32'b10011010110001100010100110110110;
		correct = 32'b10011110111111101011111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111000011110001110011100011100;
		b = 32'b11010101000011101111011110111111;
		correct = 32'b11111101011111101111011110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011010011011110111010101010;
		b = 32'b11111110110010010100011101011000;
		correct = 32'b11111111110011011110111111111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101001011111111101010101000;
		b = 32'b11011011000111000001001001111111;
		correct = 32'b11111111001111111111101011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101110111010100010111010000;
		b = 32'b01100101111101101101011000110101;
		correct = 32'b11110101111111111101011111110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000001100100101000110111001;
		b = 32'b10101111101010101110011110000001;
		correct = 32'b10101111101110101111011110111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000101001100010111010111110;
		b = 32'b01001000110110110001101000000011;
		correct = 32'b11111000111111110011111010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000001100110001111011010111;
		b = 32'b01100111110010101101101001001011;
		correct = 32'b01101111111110111101111011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010000101011111100111011100;
		b = 32'b00111011001110001100001011011100;
		correct = 32'b10111011001111011111101111011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011110110110000100100100011;
		b = 32'b11010001010000000111011111000101;
		correct = 32'b11010011110110110111111111100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010100101000111000000111111;
		b = 32'b00101010010000001100101110111001;
		correct = 32'b10101010110101001111101110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100001001101101000111000000;
		b = 32'b01000011111000101111100001101101;
		correct = 32'b11111111111001101111100111101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111000001001011101111001100;
		b = 32'b11110111000011001001010011010110;
		correct = 32'b11111111000011001011111111011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001000111011111111111111010;
		b = 32'b10100100010110011111011111001001;
		correct = 32'b10101101010111011111111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010110111001111001110110111;
		b = 32'b01101100010101010110001010110010;
		correct = 32'b11101110110111011111001110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110001111010010110010111000;
		b = 32'b01001001111101011110000011110101;
		correct = 32'b11001111111111011110110011111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010111010111100001010001001;
		b = 32'b11010000010100000111101110000011;
		correct = 32'b11111010111110111111101110001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111001011011001011000000001;
		b = 32'b00110011001000100110101101100100;
		correct = 32'b01110111001011111111111101100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110010000111001100011011100;
		b = 32'b01110111001010011101100100111010;
		correct = 32'b11110111011010111101100111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011110101110000110110110101;
		b = 32'b11101101101111000001011101001011;
		correct = 32'b11111111111111110001111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110110101111110001000111010;
		b = 32'b10010010100001010010001011111100;
		correct = 32'b10010110110101111110001011111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010010011011000010111111001;
		b = 32'b10110001000101000101000011000110;
		correct = 32'b11110011010111011101010111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011001110101000010111111011100;
		b = 32'b00101111111100001101110110011000;
		correct = 32'b00111111111101001111111111011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001100101010100100110110010;
		b = 32'b11001110011001000110111001110001;
		correct = 32'b11111111111101010110111111110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001000010010101000011000100;
		b = 32'b10000111010011000101000100100110;
		correct = 32'b11101111010011010101000111100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010111010010000011100001110;
		b = 32'b00110110110000011100001101111110;
		correct = 32'b10111110111010011100011101111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111100010100110000101000010;
		b = 32'b11100011101110101111010101100011;
		correct = 32'b11101111101110101111010101100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101110000101011111000100101;
		b = 32'b10110101101111010110000110111011;
		correct = 32'b11111101111111111111111110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011111000000000010111001110;
		b = 32'b11000000111110001100010110000101;
		correct = 32'b11001011111110001100010111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010101011110100110001101100;
		b = 32'b10000000000101110110010110011101;
		correct = 32'b11110010101111110110110111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001111000000000010101110100;
		b = 32'b10000101011000011001000000010000;
		correct = 32'b11011101111000011001010101110100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111010000010100100010100110010;
		b = 32'b00000110101011001110010101100100;
		correct = 32'b00111110101011101110010101110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010101010001010110001101011;
		b = 32'b00111011111011101100111101000000;
		correct = 32'b01111011111011101110111101101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111001100010001000101010010;
		b = 32'b10111001011010010101101011101010;
		correct = 32'b10111111011110010101101111111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100100001100101110100101111;
		b = 32'b10001101011100100100000110000110;
		correct = 32'b10001101111101100101110110101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111000011001000101100111111;
		b = 32'b11100011011111011001101101011000;
		correct = 32'b11111111011111011001101101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101010001111100110010100010;
		b = 32'b00111000110010110100011100010111;
		correct = 32'b10111101110011111100111110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111110000011101011011101100;
		b = 32'b11111100100101000000111101111011;
		correct = 32'b11111111110101011101111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000111100111011100001010010;
		b = 32'b00111001011000100010100100010100;
		correct = 32'b00111001111100111011100101010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100101000110100110011010100;
		b = 32'b11101110110110101010001101000110;
		correct = 32'b11111110111110111110111111010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110011110110101000101111100111;
		b = 32'b00001010111001010011010011010000;
		correct = 32'b10111011111111111011111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110111111011000011101010111000;
		b = 32'b11000101110111100100100111011100;
		correct = 32'b11110111111111100111101111111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101000011110110100111101110;
		b = 32'b10110100011011100111000111001100;
		correct = 32'b11111101011011110111100111101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000101101111110010101100010;
		b = 32'b01101101000000110011001111000100;
		correct = 32'b11111101101101111111011111100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000110011101111111011000101;
		b = 32'b01001010110010110100010111111001;
		correct = 32'b01011010110011111111111111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010011111011100101001001011;
		b = 32'b10110100110111000100101011001001;
		correct = 32'b11110110111111011100101011001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011011011110000111110011010;
		b = 32'b00001000001110011110000001110100;
		correct = 32'b01011011011111111110111111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101110111110011001110101001;
		b = 32'b01100001111111010010001010100000;
		correct = 32'b01111101111111110011001110101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101111000111110100111011110;
		b = 32'b00011100010111100010111110100110;
		correct = 32'b11111101111111111110111111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100000011100000001000100110;
		b = 32'b01001000100011010110001111001011;
		correct = 32'b11011100100011110110001111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101001011010000101101101100;
		b = 32'b10110001101111011001000101011001;
		correct = 32'b10111101101111011001101101111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101111111001100110110110011;
		b = 32'b01001011111101010011101110000111;
		correct = 32'b01101111111111011111111110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101110101110101011110011110;
		b = 32'b00100110011101011010000101000000;
		correct = 32'b01111111111101111111011111011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110110011100001010111000000;
		b = 32'b10001001010011011000001011101100;
		correct = 32'b10001111110011111001011111101100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000010010111011010010111111100;
		b = 32'b10110010010000011100110110000110;
		correct = 32'b11110010010111011110110111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100110110100100110001101001;
		b = 32'b00110010100011001111010001100011;
		correct = 32'b01111110110111101111110001101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110110111101101010000010011;
		b = 32'b11100011110111010101001101100011;
		correct = 32'b11101111110111111101011101110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010011000011010011001101010000;
		b = 32'b01011001010000000100000001011110;
		correct = 32'b01011011010011010111001101011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000100110010011010111000100;
		b = 32'b01111000001010011111111011101100;
		correct = 32'b01111000101110011111111111101100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101111100000011011110111010;
		b = 32'b11001010111010100101100110100001;
		correct = 32'b11011111111110100111111110111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001000000010000111001111110;
		b = 32'b10000111001000101100010010001000;
		correct = 32'b10010111001000111100111011111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011000101010001100010010011010;
		b = 32'b01010000000011000000010100111100;
		correct = 32'b01011000101011001100010110111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111001001101000110111100101;
		b = 32'b01100000010011000011010111100101;
		correct = 32'b01101111011011101011110111100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010100000100111001111001111;
		b = 32'b10110000001111000011010011111100;
		correct = 32'b11111010101111100111011111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001100011110011010100011000;
		b = 32'b00011101101101001100101100110111;
		correct = 32'b00111101101111111111111100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010001010100000000100100110;
		b = 32'b11010110010000000000101111010011;
		correct = 32'b11011110011010100000101111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011011110101000111101010011;
		b = 32'b01101001110011110110100100111000;
		correct = 32'b11101011111111111110111101111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110010101110100010110010011;
		b = 32'b11010011110001011100110111101011;
		correct = 32'b11110111110101111100110111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010100101101110111110010101;
		b = 32'b11001011011111110001110000001111;
		correct = 32'b11101011111111111111111110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000101010011101111011000101;
		b = 32'b10001100000011110010001101110001;
		correct = 32'b11001100101011111111111111110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100101100000010001000110010;
		b = 32'b00010001111011011100101011001101;
		correct = 32'b11010101111111011110101011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111110011101111100101100100011;
		b = 32'b11101000010101010100111000111111;
		correct = 32'b11111110011101111100111100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001000100111101011001011010010;
		b = 32'b01011010000101011110110000010100;
		correct = 32'b01011010100111111111111011010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010010110001000100000011001;
		b = 32'b10011010110110111100100000111101;
		correct = 32'b11011010110110111100100000111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100110111111101000110110000;
		b = 32'b10010101000010111111000110000111;
		correct = 32'b10011101110111111111000110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010011100111000111110100010;
		b = 32'b00000111111000010110001111101011;
		correct = 32'b01001111111100111110111111101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001000011000000000011111101;
		b = 32'b11010000010111010000010011000011;
		correct = 32'b11011001010111010000010011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010111001100001110011001101;
		b = 32'b10100001101111011010111111011101;
		correct = 32'b11101011111111111011111111011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110011000011001011001100001;
		b = 32'b10010100111111011111001001111110;
		correct = 32'b11110110111111011111011001111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100011011101101110111010110;
		b = 32'b10111101100001100000000100111001;
		correct = 32'b10111101111011101101110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000111011110001110111110111;
		b = 32'b00011111001001110101000101010010;
		correct = 32'b10111111111011110101110111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111111000011010001011011000;
		b = 32'b11101011110001110101110101100011;
		correct = 32'b11111111111001111111111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000100110011110001000001011;
		b = 32'b11101111001110011010100001111110;
		correct = 32'b11111111101110011110101001111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000001010111000100001110000;
		b = 32'b01110101111000010001000000001110;
		correct = 32'b11111101111010111001100001111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110100011000001011111000100101;
		b = 32'b01111011100101100110001011111011;
		correct = 32'b01111111111101101111111011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110010001000010111101010110;
		b = 32'b01100000010010101101010010000100;
		correct = 32'b01100110010011101111111111010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001001011111000001001000100;
		b = 32'b00011100001111011101010110111010;
		correct = 32'b01011101001111111101011111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010110110110001111011110110;
		b = 32'b11111101010001000111100110000100;
		correct = 32'b11111111110111110111111111110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001001100110011010011010100101;
		b = 32'b11110011101110000001001000011001;
		correct = 32'b11111011101110011011011010111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110101110001000110111001100;
		b = 32'b10101101101011010001100101111011;
		correct = 32'b11111111101111011001110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001000001010011011010000110;
		b = 32'b11100111101001110000001010000110;
		correct = 32'b11110111101001110011011010000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010111111000011000001110101;
		b = 32'b01100100010111110010011000100011;
		correct = 32'b01101110111111110011011001110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111010011110100000011100011;
		b = 32'b10100110111011101001100011001100;
		correct = 32'b11101111111011111101100011101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011100010101101101110011011;
		b = 32'b10101100000100111110110101110000;
		correct = 32'b10111111100110111111111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100011010010110010110000011110;
		b = 32'b00000010011010110010001011001101;
		correct = 32'b10100011011010110010111011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011101000101011011001111100;
		b = 32'b11101101111111010110000001100010;
		correct = 32'b11101111111111111111011001111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010100000100010010101110100;
		b = 32'b11101000001111000110110011011011;
		correct = 32'b11101010101111100110110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100100111100011011100000110;
		b = 32'b11010010010001000010110110011010;
		correct = 32'b11111110110111100011111110011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101111010001011100101111001;
		b = 32'b00111000110011111011100001000011;
		correct = 32'b11111101111011111011100101111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100100000001001001010111010;
		b = 32'b00010111000100101011111111000111;
		correct = 32'b10011111100100101011111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101010110010011110010100110;
		b = 32'b11101101000111101001100000111101;
		correct = 32'b11111101010111111011110010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110000100000011100101000100;
		b = 32'b10101001001110001101000000011100;
		correct = 32'b10101111001110001111100101011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001010010011010100100000011;
		b = 32'b11111010010000011100010010010000;
		correct = 32'b11111011010010011110110110010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100000010000000000100001110;
		b = 32'b10011100010000000101001111010000;
		correct = 32'b11011100010010000101001111011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001010001011111101000100010;
		b = 32'b01000110001001101001000100000000;
		correct = 32'b11010111011001111111101100100010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010111100001101111000100101010;
		b = 32'b00110101010110001010101100110011;
		correct = 32'b11110111110111101111101100111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110101100111111110000111010;
		b = 32'b00101111110011000001101111010011;
		correct = 32'b10101111111111111111111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000011000110100001000100011;
		b = 32'b10001001110011110100011111011101;
		correct = 32'b11001001111011110100011111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001110101011001101010110101;
		b = 32'b11000001000100011011010010110010;
		correct = 32'b11111001110101011011111010110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111110000001100011011100100;
		b = 32'b11011001101110011100001010100001;
		correct = 32'b11011111111110011100011011100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011101110011101111010001010;
		b = 32'b10100110111101110101100001101101;
		correct = 32'b10111111111111111101111011101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110000100000100010110000011;
		b = 32'b11010100110111111100110010111010;
		correct = 32'b11110110110111111100110110111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110011001000100110001110100;
		b = 32'b00010101110111110111011101001010;
		correct = 32'b10110111111111110111111101111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001011000001111110100101000;
		b = 32'b01100000010111110111110001111100;
		correct = 32'b11111001011111111111110101111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101000111011100011101011001;
		b = 32'b11101111011100011100101001101001;
		correct = 32'b11111111011111011100111101111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111111111010001011011101101;
		b = 32'b00000101000000101001000011110111;
		correct = 32'b10100111111111111001011011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111001101011011101011101000;
		b = 32'b11110010101000101001101101010000;
		correct = 32'b11111111101101111011101111111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000110111011101010000010110101;
		b = 32'b11011100010000000010000000101100;
		correct = 32'b11011110111011101010000010111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001011100110111101000011100;
		b = 32'b00010100001110101101000010100101;
		correct = 32'b01011101011110111111101010111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000110100011011010001101011000;
		b = 32'b00111011001010001100111000001000;
		correct = 32'b00111111101011011110111101011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110111101011000010101111001;
		b = 32'b10110010110100011110101011101100;
		correct = 32'b10111110111101011110111111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011100101001111110000110101;
		b = 32'b10011101100100010001000011011011;
		correct = 32'b11011111100101011111110011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111101110011111100011011010;
		b = 32'b01011100011111100111011101100111;
		correct = 32'b11111111111111111111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101100001011100001011101000;
		b = 32'b01011111110100001110001111001011;
		correct = 32'b11011111110101011110001111101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101000110101101101000100001;
		b = 32'b11110101001001011011000110001000;
		correct = 32'b11111101001111111111101110101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011111101010101111010010101;
		b = 32'b00001100101011001100010000110011;
		correct = 32'b00001111111111011101111010110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000000001100110111010010010;
		b = 32'b00011100111100001101111101100011;
		correct = 32'b11011100111101101111111111110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011101111111010000011111000011;
		b = 32'b01011001000111000110010011011101;
		correct = 32'b11011101111111010110011111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110100000110010001001011001111;
		b = 32'b00011011110010000110001100110011;
		correct = 32'b11111111110110010111001111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011011101101010011011001010;
		b = 32'b00010000101011100010000101000001;
		correct = 32'b00111011111111101010011111001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101111000010000011001111010011;
		b = 32'b11001100001011101010111100010011;
		correct = 32'b11101111001011101011111111010011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001110010001010100011111010100;
		b = 32'b10110100000110010011010101001110;
		correct = 32'b10111110010111010111011111011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111100011111001101111101111101;
		b = 32'b00100011011110100010010101110101;
		correct = 32'b00111111011111101111111101111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110101001110000011010111011;
		b = 32'b01101100100101011110001010011011;
		correct = 32'b11101110101101111110011010111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000101111111011110001000011000;
		b = 32'b01011000011110111110000000011101;
		correct = 32'b01011101111111111110001000011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000000100100001100010100110;
		b = 32'b00000100110010101011101100100100;
		correct = 32'b00010100110110101011101110100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000111110110001101101101111011;
		b = 32'b01001011011010000110010101000000;
		correct = 32'b01001111111110001111111101111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011111001011000101011001010;
		b = 32'b11000000100110010111001100011000;
		correct = 32'b11100011111111011111101111011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011010010111100011010110101;
		b = 32'b01000011100001100000000001001011;
		correct = 32'b11111011110011111100011011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100010010101100100110010110;
		b = 32'b11111100111001101101100101101111;
		correct = 32'b11111100111011101101100111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010111000001100110111000011;
		b = 32'b00000101100001100001001011000110;
		correct = 32'b00000111111001101101111111000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001100100100000001000010110;
		b = 32'b01110101110001100111111101111111;
		correct = 32'b01110101110101100111111101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001110110001001010000001111;
		b = 32'b11011101010000100111111000000111;
		correct = 32'b11111101110110101111111000001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000000000111001001110001110;
		b = 32'b11010011001101000101101000111110;
		correct = 32'b11010011001101111101101110111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001001101100011010110000000;
		b = 32'b00111111010001001000000100111110;
		correct = 32'b10111111011101101011010110111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111001000000000000110110100;
		b = 32'b10110111001010011110111011101011;
		correct = 32'b11110111001010011110111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001001001100010010011010011;
		b = 32'b01010101011011100100000000001101;
		correct = 32'b11110101011011100110010011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111111011101100011110110100;
		b = 32'b00111011001001011001011100101100;
		correct = 32'b01111111111011111101011110111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010001100110001010100000010;
		b = 32'b11010100000110010010110101000011;
		correct = 32'b11011110001110110011110101000011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110011001100101001010000011110;
		b = 32'b01011011110101000110111011010110;
		correct = 32'b11111011111101101111111011011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101101111100111001101011101;
		b = 32'b10001111011000110000011111001111;
		correct = 32'b10011111111111110111011111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101110111101010001110000100;
		b = 32'b10010011110001010100100110110111;
		correct = 32'b11011111110111111110101110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001110101001111000100110111;
		b = 32'b01001110101100100101111101100100;
		correct = 32'b01011111111101101111111101110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011110101110001110000111101;
		b = 32'b01101110110011101010101111000110;
		correct = 32'b01111111110111111011111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111111110101001011000101101;
		b = 32'b11000000011010100111001101100010;
		correct = 32'b11101111111110101111011101101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100110000110100011110110010100;
		b = 32'b11111100110101010110101111000001;
		correct = 32'b11111110110111110111111111010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100000101000001111001001011;
		b = 32'b01101101001110010101000100010010;
		correct = 32'b01101101001111010101111101011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100100110100011100010100101;
		b = 32'b11000111011010101010001000100001;
		correct = 32'b11110111111110101011101010100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000100111011001000101011010001;
		b = 32'b00101000111110111001001011110000;
		correct = 32'b00101100111111111001101011110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110010000100100100111111010111;
		b = 32'b11110110101100001100001001001010;
		correct = 32'b11110110101100101100111111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011100010010100101011001110;
		b = 32'b11111011110111111101010010010101;
		correct = 32'b11111011110111111101111011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001100010001111000011001100;
		b = 32'b10101110010100010010010000011101;
		correct = 32'b10111111110110011111010011011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110100100101101111101110100;
		b = 32'b00001101101011111100101111110111;
		correct = 32'b00011111101111111101111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011010110100101111001001000111;
		b = 32'b00001101111100001101001100010001;
		correct = 32'b11011111111100101111001101010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011101101010110000111101011;
		b = 32'b00001101110110011110000100010011;
		correct = 32'b01001111111111011110000111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000110101000110001000000010;
		b = 32'b01111001011011100100010100011101;
		correct = 32'b11111001111111100110011100011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110001011110001011010001110011;
		b = 32'b10001001101000011110101011111000;
		correct = 32'b10111001111110011111111011111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011111011001011111011111111;
		b = 32'b00000010101110000010011101111011;
		correct = 32'b00110011111111001011111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111001011000001111100011011101;
		b = 32'b10011000111010111100011010011101;
		correct = 32'b10111001111010111111111011011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111001000110101010011001001;
		b = 32'b00000100000001101100011100101000;
		correct = 32'b00001111001001111101011111101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100110001100101001010011000;
		b = 32'b01100001001110000101001101101011;
		correct = 32'b01101101111111100101001111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010111010111111001111000110;
		b = 32'b10000011110101100101111001001010;
		correct = 32'b11101011111111111111111111001110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000101111011100011111100010;
		b = 32'b01101001101100111010010110110111;
		correct = 32'b01111001101111111110011111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000001010010111001101011110;
		b = 32'b10100111001010111000110101111111;
		correct = 32'b11100111001010111111111101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110111101001101001010001001100;
		b = 32'b00100010010011100011100111110110;
		correct = 32'b11110111111011101011110111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001010010110010011011010010;
		b = 32'b11110010111101011000111001110010;
		correct = 32'b11111011111111111010111011110010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101000101111010001100001100010;
		b = 32'b00100101011111010111010100101010;
		correct = 32'b01101101111111010111110101101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001010110110010011110011100;
		b = 32'b10010010010101111010000111001101;
		correct = 32'b11010011010111111010011111011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100111110000011010111001011000;
		b = 32'b10000001000100111001100000010001;
		correct = 32'b11100111110100111011111001011001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011001001110010100011010111;
		b = 32'b11100111001011110100101001010101;
		correct = 32'b11111111001011110110101011010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001010110000011010001000010;
		b = 32'b01100001001110010101001000001100;
		correct = 32'b01101001011110010111011001001110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110011011110100101101000100;
		b = 32'b11100000101010001000111101100101;
		correct = 32'b11110110111011111100111101100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011100000000011100000111110;
		b = 32'b10110000001111110011100000011101;
		correct = 32'b11111011101111110011100000111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111111010101111111111100101;
		b = 32'b10010111111100111111001001011001;
		correct = 32'b11011111111110111111111111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101101101100110011101110010;
		b = 32'b01101100111001011101010011110000;
		correct = 32'b11111101111101111111011111110010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011011100000010100101110111000;
		b = 32'b10010111010101001100000000010101;
		correct = 32'b11011111110101011100101110111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111110010010001000100011111101;
		b = 32'b11011010100000011110001111100101;
		correct = 32'b11111110110010011110101111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011000011100011000000010100;
		b = 32'b00000110010000000100101101101000;
		correct = 32'b10001111010011100111101101111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100110001100111000101101001;
		b = 32'b11100101011001110000010001000110;
		correct = 32'b11111101111001110111010101101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110011011111111011001000110;
		b = 32'b00010101111100110010111011000011;
		correct = 32'b00111111111111111111111011000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011001110010001101110010010;
		b = 32'b00001100001101010100111110011111;
		correct = 32'b01111111001111010101111110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001101111100110011100100101;
		b = 32'b11101100001001100100101011100010;
		correct = 32'b11101101101111100110111111100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110010001100010101010101001;
		b = 32'b10110011100000001010000110101101;
		correct = 32'b10110111110001101010101110101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011011010011011000000100110;
		b = 32'b11011001101111110100100001001111;
		correct = 32'b11111011111111111111100001101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000111000100010010010110011;
		b = 32'b00110111100101000011010001001001;
		correct = 32'b10110111111101100011010011111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001100000010010001000101011;
		b = 32'b00110100010101100000000000111000;
		correct = 32'b11111101110101110010001000111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000101010001001111011101110;
		b = 32'b01010010111000011010011010100000;
		correct = 32'b11010010111010011011111011101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100010000001000110100011110000;
		b = 32'b11001110001011000101101010010010;
		correct = 32'b11101110001011000111101011110010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101000101000001010111101100;
		b = 32'b01000010011100000110111010110111;
		correct = 32'b01000111011101000111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111111000101000001111110011;
		b = 32'b00100000001110001111000011110100;
		correct = 32'b11111111111110101111001111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111100010000011110010110110;
		b = 32'b01101100001101011100101100011000;
		correct = 32'b01101111101111011111111110111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010100000000100101100100110;
		b = 32'b00101000011011010011000010010011;
		correct = 32'b00111010111011010111101110110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000110101001011011110010000;
		b = 32'b11000011110101110011110011101011;
		correct = 32'b11011011110101111011111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101101101010111001010100011;
		b = 32'b01000010110100110100010110111101;
		correct = 32'b01010111111101110111011110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011011011110011011011110010;
		b = 32'b11101001010111101001001101010101;
		correct = 32'b11111011011111111011011111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111011110110111110011001000;
		b = 32'b01100011111010100101000001110100;
		correct = 32'b11100111111110110111110011111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111000111000001110100001000000;
		b = 32'b11100101011111101000110110110100;
		correct = 32'b11111101111111101110110111110100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100110101101010011011111110;
		b = 32'b11010101111101001001010001111000;
		correct = 32'b11010101111101101011011011111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001101010010100100101000110;
		b = 32'b11111010110011010100110100100110;
		correct = 32'b11111011111011010100110101100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000110111010000110111010000;
		b = 32'b10101101110100011010110110001111;
		correct = 32'b10111101110111011010110111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010001011001110101111101111;
		b = 32'b10110001101100100111111010001110;
		correct = 32'b10111011101111101111111111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011110111100111000101101010;
		b = 32'b10001111011010111111000011111111;
		correct = 32'b10001111111111111111000111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101111011101011010011000110;
		b = 32'b10100110101010011111000111011100;
		correct = 32'b10101111111011111111010111011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001101010111111010001010011;
		b = 32'b00001010011000110010110101101100;
		correct = 32'b01011011111010111111110101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001001111101000111000011011;
		b = 32'b00001010001000110111111111110101;
		correct = 32'b10101011001111111111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000000101111000100100100100100;
		b = 32'b01110000101100001010011011000101;
		correct = 32'b11110000101111001110111111100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100111000110010000111011000;
		b = 32'b10000111010111110001100010011100;
		correct = 32'b10001111111111110011100111011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101111000100110100000111101;
		b = 32'b10111111011110111001110011011111;
		correct = 32'b11111111111110111111110011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001100011110100010011101001;
		b = 32'b00011000010010110011110101010101;
		correct = 32'b11011001110011110111110111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111101010010000011000100100;
		b = 32'b10100110100010100100100100011111;
		correct = 32'b11110111101010110100111100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010111100101000110111101110;
		b = 32'b01001000101100101011011110100100;
		correct = 32'b11001010111100101011111111101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110001101100110001101110101101;
		b = 32'b10101001100000101110001101011110;
		correct = 32'b11111001101100111111101111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100011101100000001111010011;
		b = 32'b01000101100010001001010000101001;
		correct = 32'b11111101111111101001011111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101101010011000110011010011;
		b = 32'b00010110110010100000010110111111;
		correct = 32'b10111111111010111000110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111001001111010110111011100;
		b = 32'b00100011010110110010000110010011;
		correct = 32'b00101111011111111010110111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000100100010101101010110001100;
		b = 32'b01000100111101010100010101010100;
		correct = 32'b11000100111111111101010111011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000011001100011110100110111;
		b = 32'b00000011001010110001011011101101;
		correct = 32'b10011011011011110011111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101100001100100111100100110;
		b = 32'b11110001000010010001010110011010;
		correct = 32'b11111101100011110101111110111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000000101001110110110101010;
		b = 32'b00000100100011000110001110110101;
		correct = 32'b00010100100111001110111110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010111011100000110010100100;
		b = 32'b01000000001110100000010001000001;
		correct = 32'b01101010111111100000110011100101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001110010010101001101011011;
		b = 32'b00001011110000011010110100010101;
		correct = 32'b01101011110010011111111101011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110011000111111010010011010;
		b = 32'b00100010011110110101101001111101;
		correct = 32'b01111110011110111111111011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011110000101110000100100010001;
		b = 32'b01010110101100011001001101001101;
		correct = 32'b01011110101101111001101101011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000110110000001101100000100;
		b = 32'b10001110010110001011101001001000;
		correct = 32'b11001110110110001011101101001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011010010101101001001111110;
		b = 32'b10101010011111011000101101001100;
		correct = 32'b11101011011111111101101101111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101111111010101100001110010;
		b = 32'b01011000110110001000010101011010;
		correct = 32'b01011101111111011101110101111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111110111101110011010111100001;
		b = 32'b11001101100111011100101111101000;
		correct = 32'b11111111111111111111111111101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001111010111110100100101111;
		b = 32'b01111110100111101011011111010010;
		correct = 32'b11111111111111111111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001110100011001001000100011;
		b = 32'b11001101111101010001101011001010;
		correct = 32'b11101101111101011001101011101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001100111101101111110000111;
		b = 32'b10011001111101011101001111000110;
		correct = 32'b11011001111111111101111111000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110101001011011000101111000;
		b = 32'b00101110010100111010010100001001;
		correct = 32'b10111110111101111011010101111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110110100010001010000101000;
		b = 32'b11011101101000001101110100001100;
		correct = 32'b11111111111100011101110100101100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110111010001111010101100001100;
		b = 32'b10100110111010000111111010111001;
		correct = 32'b10110111111011111111111110111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011000011010111101010100111000;
		b = 32'b00101100001101000010000001000000;
		correct = 32'b11111100011111111111010101111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001001001011101011000100001;
		b = 32'b11001000111111011110001101001010;
		correct = 32'b11011001111111011111011101101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100110100111101101011101011100;
		b = 32'b11011011000001101111010000100001;
		correct = 32'b11111111100111101111011101111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111000111011010111110101010;
		b = 32'b01001011010011101101010100100110;
		correct = 32'b11011111010111111111111110101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000010011100011000010101000;
		b = 32'b11010110100100100011010000101011;
		correct = 32'b11011110110111100011010010101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010010111000011010110010100011;
		b = 32'b11010110001100000101011111110110;
		correct = 32'b11010110111100011111111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110001101101111000110000001111;
		b = 32'b01001011100111010000110111101101;
		correct = 32'b01111011101111111000110111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010111101100011011110101010;
		b = 32'b10000011011010000101010010000001;
		correct = 32'b10111011111111100111011110101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010011010000011110001011111;
		b = 32'b01111101101111110001100011010101;
		correct = 32'b01111111111111110011110011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110010000100000001011001000110;
		b = 32'b10101110010001011001110000111011;
		correct = 32'b10111110010101011001111001111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001110111111111010100100001;
		b = 32'b10001011101100101101010111110011;
		correct = 32'b10101011111111111111010111110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010000011111010101110100000000;
		b = 32'b10111010001000100010110010010101;
		correct = 32'b11111010011111110111110110010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000110101110101110010001101;
		b = 32'b10001101100100111000010101001101;
		correct = 32'b11011101110101111101110111001101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001100000000000100110010110;
		b = 32'b11000001101101100001100101010110;
		correct = 32'b11000001101101100001100111010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100111000111100100110101011;
		b = 32'b11111100101011011101011000011100;
		correct = 32'b11111100111011111101111110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010101110011000100011010000;
		b = 32'b01111101010110011100010100000110;
		correct = 32'b01111111111110011100110111010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000111001000100110110001000011;
		b = 32'b11111110110011110010000110101011;
		correct = 32'b11111111111011110110110111101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110111010000001011011101001;
		b = 32'b10100101010001001001000100111011;
		correct = 32'b11110111111011001001011111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011011100101000011110000111;
		b = 32'b10000000101110101101000001101110;
		correct = 32'b10111011111110101101011111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111101101111111111100100001;
		b = 32'b00011111001010111110101100001111;
		correct = 32'b01011111101111111111111100101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010100101001010010011100100001;
		b = 32'b01101000100011011100110110000001;
		correct = 32'b01111100101011011110111110100001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111111110111101110110100011111;
		b = 32'b01111000011010000001011110101001;
		correct = 32'b11111111111111101111111110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110110100000100000101001011;
		b = 32'b00111101100000110000010011001110;
		correct = 32'b11111111110100110100010111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010001110001100000010001111;
		b = 32'b01010000101000011100001010111001;
		correct = 32'b11110010101110011100001010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011101101010000110111010110011;
		b = 32'b10001010010100000001100010110100;
		correct = 32'b10011111111110000111111010110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011101011110010101000101100;
		b = 32'b01010100011001010010101110010110;
		correct = 32'b11110111111011110010101110111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001010000111111110111010001100;
		b = 32'b10010111001010001011011011011111;
		correct = 32'b11011111001111111111111011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010110100110100011001001110;
		b = 32'b10110011101000110110110000100111;
		correct = 32'b11110011111100110110111001101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010001011111101010011010000100;
		b = 32'b01010010111010111111110101010011;
		correct = 32'b01010011111111111111111111010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110011010000000011010110101;
		b = 32'b00000000000111001100110000011100;
		correct = 32'b01001110011111001100111010111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001111010010110100010100011;
		b = 32'b10110110010001001010011110000001;
		correct = 32'b10111111111011011110111110100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010001101110100000010000110;
		b = 32'b01000001100010110110000011010010;
		correct = 32'b11000011101111110110000011010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001101010110000111101101001;
		b = 32'b11111101011100100111001110101010;
		correct = 32'b11111101111110110111111111101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010010110011101101100111110;
		b = 32'b01101100010001011000010001101000;
		correct = 32'b01101110010111011101111101111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110011001100100011110001100110;
		b = 32'b00101110111010001100111001110000;
		correct = 32'b01111111111110101111111001110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011001111100101010101001100000;
		b = 32'b01101011010010001000110010110011;
		correct = 32'b01111011111110101010111011110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001000101001110101101010001;
		b = 32'b01000000011101010000110110111101;
		correct = 32'b11001001011101011110111111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001101101000001011000101000;
		b = 32'b01001011110001100011010100001001;
		correct = 32'b11011011111101100011011100101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111101011111100000000011100;
		b = 32'b10000110100101010011100010100111;
		correct = 32'b10010111101111111111100010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101111100101110010111101001;
		b = 32'b10000110101111000100110111001100;
		correct = 32'b10010111111111101110110111101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000110001101100011010001111;
		b = 32'b00111101011000111111001100010100;
		correct = 32'b00111101111001111111011110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000010000001011001001001101;
		b = 32'b10010000011010101100100000001100;
		correct = 32'b10110000011010101111101001001101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100110000110101011010011111;
		b = 32'b10011000010110111101100100001101;
		correct = 32'b11011100110110111101111110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000101010000101101101010001;
		b = 32'b11000001111010101000001100110011;
		correct = 32'b11100001111010101101101101110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110110000100100111010011011111;
		b = 32'b10110000001001111110000100100100;
		correct = 32'b10110110001101111111010111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110110110100001011110001010;
		b = 32'b01000011100100001000000101001110;
		correct = 32'b11001111110110101001011111001110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100111010100001011110011011011;
		b = 32'b00010100101001110010100110010001;
		correct = 32'b10110111111101111011110111011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010000011101000010000000010;
		b = 32'b01100001011111011001101000001111;
		correct = 32'b01100011011111111001111000001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110011011001010001110110100;
		b = 32'b01110001111111011101110000001011;
		correct = 32'b11111111111111011111111110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101111101101001111001101001;
		b = 32'b00111111111011100110000110011000;
		correct = 32'b11111111111111101111111111111001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010001100111001000100010110;
		b = 32'b10100001010011011001101011110000;
		correct = 32'b10111011011111111001101111110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111101010000101001010110111;
		b = 32'b11111011100101111010110000101110;
		correct = 32'b11111111101111111111111010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011000111010111001111100110;
		b = 32'b01001001011000100100001100101011;
		correct = 32'b01001011011111110111001111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010000011010001100110101111111;
		b = 32'b01011101100100010011100000101011;
		correct = 32'b11011101111110011111110101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100101000110100000110001000001;
		b = 32'b10100100110110101110100111100111;
		correct = 32'b10100101110110101110110111100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010101010110000001000101000;
		b = 32'b01111001100001100101110110101000;
		correct = 32'b01111011101011110101111110101000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111000001000001011111111100;
		b = 32'b01101110010111101111110001001000;
		correct = 32'b01111111010111101111111111111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000010100101100100001110011001;
		b = 32'b11110010100000101110001010111010;
		correct = 32'b11110010100101101110001110111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110000111000010000101101110;
		b = 32'b10101011000110001111100110100000;
		correct = 32'b11101111000111001111100111101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100010000010000111000110110;
		b = 32'b10110111110101100001111110011111;
		correct = 32'b11111111110101110001111110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011010000010001100110111011001;
		b = 32'b01010100011011110000100110011010;
		correct = 32'b11011110011011111100110111011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011011001000000100100111111111;
		b = 32'b10100110101010001000110111011011;
		correct = 32'b11111111101010001100110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010011101010110111000001010;
		b = 32'b00101001110010000000000010111001;
		correct = 32'b00101011111111010110111010111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111111111100101011001000010101;
		b = 32'b01110010110001111101001100010101;
		correct = 32'b11111111111101111111001100010101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011000101110100110111001100;
		b = 32'b00100011000011110110111101000100;
		correct = 32'b10111011000111110110111111001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111100100101011110001101101;
		b = 32'b11000001100111101101101110101000;
		correct = 32'b11010111100111101111111111101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101101010011000101110111111010;
		b = 32'b00111000110100100110000000100111;
		correct = 32'b10111101110111100111110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000101100100011011000100111000;
		b = 32'b11010100010011111011000001001101;
		correct = 32'b11010101110111111011000101111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100111100111000010001001011;
		b = 32'b01001011111000100100110001110011;
		correct = 32'b01111111111100111100110001111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101010111111111110001110110;
		b = 32'b11100100101001001010100100100011;
		correct = 32'b11100101111111111111110101110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010101011010101111101100110;
		b = 32'b01111101100111110011110100000110;
		correct = 32'b11111111101111110111111101100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011101011001001111101000010;
		b = 32'b11101001110011111100010011000100;
		correct = 32'b11111011111011111101111111000110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100001010000001111100111001101;
		b = 32'b10010011110101001101000110001010;
		correct = 32'b10110011110101001111100111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100100101100000110010011111;
		b = 32'b01111011000110010001110110010010;
		correct = 32'b11111111100111110001110110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101111011000011100010000111;
		b = 32'b10010110110100010010000100010110;
		correct = 32'b11011111111111010011100110010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100000001110111100110100011111;
		b = 32'b01100011000110110000101000110100;
		correct = 32'b01100011001110111100111100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011101000001001001011100011010;
		b = 32'b00101011010100011011010100001001;
		correct = 32'b10111111010101011011011100011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010011000010110000011111101001;
		b = 32'b10011010100101000101110011000100;
		correct = 32'b10011011100111110101111111101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110001111101100011110010111011;
		b = 32'b00011010000100001000111100101100;
		correct = 32'b10111011111101101011111110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001000110011010110100101110010;
		b = 32'b01010111110010111000111001111000;
		correct = 32'b01011111110011111110111101111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010111101111111110001000011110;
		b = 32'b00001111000010000110111010101001;
		correct = 32'b01011111101111111110111010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100110000000110100101010101000;
		b = 32'b11010100110110000010001001111100;
		correct = 32'b11110110110110110110101011111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000011000110000000100101001100;
		b = 32'b00011100101100101011010100010001;
		correct = 32'b10011111101110101011110101011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101100111110000011011001011011;
		b = 32'b10011010111010100010011111011000;
		correct = 32'b11111110111110100011011111011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100100100011111101110010100;
		b = 32'b01100011001100101010100100001000;
		correct = 32'b01110111101100111111101110011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101011101000001101000101011;
		b = 32'b10101111111011010011011011011100;
		correct = 32'b10111111111111010011111011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100000101110000101001110011;
		b = 32'b01110101011010011011000000011100;
		correct = 32'b11111101011111111011101001111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001100010110000011000101101100;
		b = 32'b10111110100010111011001101000111;
		correct = 32'b10111110110110111011001101101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111011001110010111011110010100;
		b = 32'b00010100101000100000001011101100;
		correct = 32'b00111111101110110111011111111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100001100000110100000000000000;
		b = 32'b00011101111001011000001010000010;
		correct = 32'b01111101111001111100001010000010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110111001011010100011001100;
		b = 32'b11100101001110101101100010001000;
		correct = 32'b11101111111111111111100011001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101111011000001100110001000;
		b = 32'b11101100000011001111001111101001;
		correct = 32'b11101101111011001111101111101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001000011010101100011000000;
		b = 32'b01001111100110011010101111101011;
		correct = 32'b01001111100111011111101111101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001100011000101111101011011;
		b = 32'b00010110111000000101100111011011;
		correct = 32'b10111111111011000101111111011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101011011111100001100101111100;
		b = 32'b10010110110111010101111110111011;
		correct = 32'b11111111111111110101111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001110100000101110100000101010;
		b = 32'b10001100110111101111001001110011;
		correct = 32'b11001110110111101111101001111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010010000001001101001110000010;
		b = 32'b11110001010011001011010000101111;
		correct = 32'b11110011010011001111011110101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000100111001111110101010100;
		b = 32'b01010001001000001100100110101100;
		correct = 32'b01110001101111001111110111111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101001001110010010000000010011;
		b = 32'b00110001011100100111100000111100;
		correct = 32'b01111001011110110111100000111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011100000110000110110011011;
		b = 32'b00010100010001010101101011010110;
		correct = 32'b11011111110001110101111111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101001111010100011010100111;
		b = 32'b01100011000010001100101010000010;
		correct = 32'b11100111001111011100111010100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011110011101010110000100101100;
		b = 32'b00010101100001000101111110101100;
		correct = 32'b11011111111101010111111110101100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100110111010111111110100000001;
		b = 32'b01110101000110001111100100011100;
		correct = 32'b11110111111110111111110100011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011111001001011001111110101;
		b = 32'b10010101110111001010111001110010;
		correct = 32'b11010111111111001011111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101110001100001101011100011000;
		b = 32'b00010110101000101001111101110100;
		correct = 32'b00111110101100101101111101111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101000011001010001000001011;
		b = 32'b11111110001000101100110000001011;
		correct = 32'b11111111001011101110111000001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010110101111011011001110110;
		b = 32'b11100110011001011100010101110010;
		correct = 32'b11100110111101111111011101110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110001100100100100011101100;
		b = 32'b00001010100000001101000101000010;
		correct = 32'b10011110101100101101100111101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010111100100010001111111000;
		b = 32'b00001000100000001000110110111111;
		correct = 32'b10111010111100101010111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100100111111010110111100100;
		b = 32'b11010001001100001011111011001101;
		correct = 32'b11011101101111111011111111101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00100000111010001100100100010100;
		b = 32'b00101010100110110011110001100001;
		correct = 32'b00101010111110111111110101110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010100110111011111110010000;
		b = 32'b11000110111111000110001100001101;
		correct = 32'b11101110111111111111111110011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110100100100110001010000010;
		b = 32'b11110011011110000000011010110001;
		correct = 32'b11110111111110100110011010110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110010001011001011111110111;
		b = 32'b11110010010100000000001111011100;
		correct = 32'b11111110010101011001011111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000001101110111010100111111;
		b = 32'b00110010100111111100010001100110;
		correct = 32'b01110010101111111111010101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011100111010001101000101111;
		b = 32'b00100111000110011010000110011011;
		correct = 32'b10111111100111011011101110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101000100101110100000001101010;
		b = 32'b11110101001001010111011011110111;
		correct = 32'b11111101101101110111011011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001011110011111111110100011110;
		b = 32'b01000101010001111001100101110001;
		correct = 32'b11001111110011111111110101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010011010110001111010101000;
		b = 32'b00010100001001000001001011000001;
		correct = 32'b00111110011011110001111011101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011100000101100011001100101101;
		b = 32'b01111001010010001101110101010110;
		correct = 32'b01111101010111101111111101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011011001010011111000111111101;
		b = 32'b01011111111001111011001001011011;
		correct = 32'b11011111111011111111001111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010111010101011001000010100000;
		b = 32'b10100100110110110011111000001010;
		correct = 32'b10110111110111111011111010101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001101110010110000110000011110;
		b = 32'b11100001010011101010000011100100;
		correct = 32'b11101101110011111010110011111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100011100011111100111100001011;
		b = 32'b01110100011101111001110000100100;
		correct = 32'b01110111111111111101111100101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110111101101010111011000010;
		b = 32'b10000111000011101010101101000111;
		correct = 32'b11010111111111101010111111000111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001011111000000010111000001;
		b = 32'b01001000001111011000111110111110;
		correct = 32'b01001001011111011000111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011100111101010101111011011010;
		b = 32'b10101011001010110010110100000100;
		correct = 32'b10111111111111110111111111011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000111011111000000010001011110;
		b = 32'b00101100011010101101000101101010;
		correct = 32'b11101111011111101101010101111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011100010010110111111010001;
		b = 32'b00100100111000011100100010010000;
		correct = 32'b00101111111010011110111111010001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001010011110001100101001101110;
		b = 32'b00110011111001011101100101100011;
		correct = 32'b11111011111111011101101101101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001100000010111001110100001100;
		b = 32'b11001110010001111010001110011101;
		correct = 32'b11001110010011111011111110011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001001100000100001010000111000;
		b = 32'b01110100111100001101101100010000;
		correct = 32'b01111101111100101101111100111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111110010111010010101000100111;
		b = 32'b11111010101011100011000000011010;
		correct = 32'b11111110111111110011101000111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110100000100000100011000100101;
		b = 32'b11111100100101101010101010110010;
		correct = 32'b11111100100101101110111010110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110011000000000011010010010;
		b = 32'b10110010111000001111000011010110;
		correct = 32'b10111110111000001111011011010110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101000010011111111101011000101;
		b = 32'b00000001001000001101001100110100;
		correct = 32'b11101001011011111111101111110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101000111111001110011100100;
		b = 32'b01000110110011111101011100101010;
		correct = 32'b11111111110111111101111111101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111001111111011001101111111;
		b = 32'b11000011001110000110001011101001;
		correct = 32'b11001111001111111111001111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111100110111011011101111111;
		b = 32'b10101000101100100111011011100100;
		correct = 32'b11101111101110111111011111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000010010110000110100001111;
		b = 32'b00101011111010010010000100101110;
		correct = 32'b10111011111010110010110100101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001110011011101000010111010;
		b = 32'b01000011000100010000011100000100;
		correct = 32'b11010011110111011101011110111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101000001000000100011010000110;
		b = 32'b01111000000100011111000001011000;
		correct = 32'b11111000001100011111011011011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000001010101000010111000111001;
		b = 32'b11100111010000010001000100110101;
		correct = 32'b11100111010101010011111100111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110000000000000011010111001;
		b = 32'b00011010001101111110111101001011;
		correct = 32'b11011110001101111110111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00111111111110000001000000100111;
		b = 32'b01001000010100111000000110001001;
		correct = 32'b01111111111110111001000110101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101110100100001111011001111110;
		b = 32'b10100100010111110001100000101110;
		correct = 32'b10101110110111111111111001111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100011011110000111111111101;
		b = 32'b10111001011011110110010001001111;
		correct = 32'b11111101011011110110111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111000110110011011101011111;
		b = 32'b00101000100101100100011010101001;
		correct = 32'b11101111100111110111011111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001101001100100010000011100011;
		b = 32'b00100001001111000101110110110101;
		correct = 32'b11101101001111100111110111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100100001011110001000011100111;
		b = 32'b11101001110011100110110111110111;
		correct = 32'b11101101111011110111110111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010011100101110100001110101;
		b = 32'b10110111110100111100100111100111;
		correct = 32'b10111111111100111110100111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110010110100010101101111011101;
		b = 32'b10000001110000111111001101110011;
		correct = 32'b10110011110100111111101111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101001010101111001101110011;
		b = 32'b11010110111101111110100111110110;
		correct = 32'b11010111111111111111101111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011000001101111001010010101000;
		b = 32'b00101010000100100001101111010000;
		correct = 32'b01111010001101111001111111111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100010000101100111001001001011;
		b = 32'b00111010101100011010100001111111;
		correct = 32'b01111010101101111111101001111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011111011010010001111111010110;
		b = 32'b10000001101100010010010010101010;
		correct = 32'b11011111111110010011111111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000011010110110000110010101110;
		b = 32'b11011000001011001011111111010001;
		correct = 32'b11011011011111111011111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101110001100101100111001010;
		b = 32'b10001111001011100001101000100001;
		correct = 32'b11011111111011100101101111101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101001111101010111101001011000;
		b = 32'b10011000101001000100001111111111;
		correct = 32'b10111001111101010111101111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101100110000101000010111011;
		b = 32'b00100110010111101011010101111101;
		correct = 32'b10110111110111101111010111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110000011111101100110100001;
		b = 32'b01010001001111110111000101010110;
		correct = 32'b11011111001111111111100111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011111111111001011111010100;
		b = 32'b11000100100110100110011110111100;
		correct = 32'b11000111111111111111011111111100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011010000010000000010011110;
		b = 32'b11010111111000100010101110001010;
		correct = 32'b11111111111000110010101110011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010000011101110000000001011;
		b = 32'b01010011111000000001000101100001;
		correct = 32'b11111011111011101111000101101011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001110001010111000110010101110;
		b = 32'b11001110110000111100001101001110;
		correct = 32'b11001110111010111100111111101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111010001110110100011101100110;
		b = 32'b10110101110010000110000000000011;
		correct = 32'b11111111111110110110011101100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001100011011110001000011100;
		b = 32'b10110100111011001011010110011111;
		correct = 32'b10111101111011011111011110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010110011010001011110001101;
		b = 32'b00101100100100011110010100100111;
		correct = 32'b10101110110111011111011110101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100100101010011000010000111010;
		b = 32'b11100001101011100001000001011000;
		correct = 32'b11100101101011111001010001111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001111001010111010010001101;
		b = 32'b10001011001111100000110110010010;
		correct = 32'b11101011111111110111110110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010011001000110111111111110111;
		b = 32'b11000100000011101110111111010111;
		correct = 32'b11010111001011111111111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000100100110000011001000111100;
		b = 32'b00001101000100010001000110101011;
		correct = 32'b01001101100110010011001110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110011000110001101010111000000;
		b = 32'b10100000000110100001011110010000;
		correct = 32'b10110011000110101101011111010000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000010011010101001001111101;
		b = 32'b01111001000110111000011110111000;
		correct = 32'b11111001010111111101011111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010111110100111000001001101;
		b = 32'b00010010001010110010000010111111;
		correct = 32'b00011010111110110111000011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000110110010101011100011110;
		b = 32'b10001101100010001100001100101000;
		correct = 32'b10011101110110011101011100111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010101110011101110010011101111;
		b = 32'b01101100000000000110110010001001;
		correct = 32'b11111101110011101110110011101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110000100011011101100100110101;
		b = 32'b11001110010101011011101001011111;
		correct = 32'b11111110110111011111101101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001010100000101000111010000000;
		b = 32'b00010000011101110101110010100110;
		correct = 32'b00011010111101111101111010100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011010010010001111111110101;
		b = 32'b01001101000001110110101000101011;
		correct = 32'b11101111010011110111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101111001011101101100001011110;
		b = 32'b00011110000011010001100100100000;
		correct = 32'b00111111001011111101100101111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110001001010011010010001001;
		b = 32'b01010111011101011010110100010010;
		correct = 32'b11010111011101011011110110011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011000011011100101010111101;
		b = 32'b00011111101011000010111101000101;
		correct = 32'b01111111101011011110111111111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010111100111101111010100111110;
		b = 32'b11010011000111011001111000000011;
		correct = 32'b11010111100111111111111100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001101110100110011010000001110;
		b = 32'b00011001100110001111100101010100;
		correct = 32'b01011101110110111111110101011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111100111010010001111100101;
		b = 32'b10000000010000010011110111000011;
		correct = 32'b10011111110111010011111111100111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110000011011100111101010110011;
		b = 32'b01111001101101011000000111110111;
		correct = 32'b01111001111111111111101111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010110110101000010010011110100;
		b = 32'b01011100111011101101000101111010;
		correct = 32'b01011110111111101111010111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111011100110101011111111101100;
		b = 32'b01100110010100000011110011100111;
		correct = 32'b11111111110110101011111111101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001111110100000001001101100011;
		b = 32'b11111110110000001100110110000011;
		correct = 32'b11111111110100001101111111100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011010111101000110111101111111;
		b = 32'b00010010111010101010101000001011;
		correct = 32'b00011010111111101110111101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001000101010001011000100111110;
		b = 32'b10111101001001001000011000001011;
		correct = 32'b11111101101011001011011100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111010100101011111000011010010;
		b = 32'b11010011101010110100000011011000;
		correct = 32'b11111011101111111111000011011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001111110001001000101100010010;
		b = 32'b01011011010111110101011100010010;
		correct = 32'b01011111110111111101111100010010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111101011000100110010110111111;
		b = 32'b10110000011000011011001111110000;
		correct = 32'b10111101011000111111011111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100010100001010000011111000;
		b = 32'b00100101110100111001010110100000;
		correct = 32'b11101101110100111011010111111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000100110001110100101110001000;
		b = 32'b01011110010000010010100000011000;
		correct = 32'b11011110110001110110101110011000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011011101000011011000001100011;
		b = 32'b10000101010000100111000101100010;
		correct = 32'b10011111111000111111000101100011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111101011011111100000011010;
		b = 32'b11101011111011100001010111000101;
		correct = 32'b11101111111011111111110111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00110000110000111000111001010010;
		b = 32'b00110010001101001010101010011001;
		correct = 32'b00110010111101111010111011011011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001111100001101001001010111;
		b = 32'b11100011100000011010111101100010;
		correct = 32'b11111011111100011111111101110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000011110111001100001000000111;
		b = 32'b00011110001110110111000110010100;
		correct = 32'b00011111111111111111001110010111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001001101011111011010011110000;
		b = 32'b10000110000101001111000110010110;
		correct = 32'b10001111101111111111010111110110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111101001110000100000101110100;
		b = 32'b11010011000111101001100101100011;
		correct = 32'b11111111001111101101100101110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111100101100001001011001100001;
		b = 32'b00111110000100110110000101110001;
		correct = 32'b10111110101100111111011101110001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110110110111001011101000010000;
		b = 32'b10100111100000111001011010111010;
		correct = 32'b10110111110111111011111010111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011000100000000111001000110010;
		b = 32'b10001011010111010100111101010101;
		correct = 32'b10011011110111010111111101110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011001010011001000111110101100;
		b = 32'b00100010010011111000000100111011;
		correct = 32'b10111011010011111000111110111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010001110011001110110110011101;
		b = 32'b00011101000000110001001111111110;
		correct = 32'b10011101110011111111111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011111111001011111110101000;
		b = 32'b01110000000000011100110010111010;
		correct = 32'b11111011111111011111111110111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001111010010111001111001000;
		b = 32'b01110100110100010100011001110010;
		correct = 32'b01111101111110010111011111111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101010110100010111001101110010;
		b = 32'b11101000011111100110110101001100;
		correct = 32'b11101010111111110111111101111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100010000000011010001000010000;
		b = 32'b11011010001001001000001100011101;
		correct = 32'b11111010001001011010001100011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000000101011000010000101011011;
		b = 32'b10101101101000000100100110111110;
		correct = 32'b10101101101011000110100111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010001010111001001001010011;
		b = 32'b11011001000110000100001000111010;
		correct = 32'b11111011001110111101001001111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101010011100011111101000110011;
		b = 32'b01100110011000000101011010001101;
		correct = 32'b01101110011100011111111010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110000101101001111100100100;
		b = 32'b00001111100100111011111111100110;
		correct = 32'b11101111100101111011111111100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01110010110010110010101011010101;
		b = 32'b01000100011101111010110101100000;
		correct = 32'b01110110111111111010111111110101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001001100101010101100100100001;
		b = 32'b00111010000011111000000001010010;
		correct = 32'b00111011100111111101100101110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100011010011100111110010011011;
		b = 32'b10110111011010110011001011101001;
		correct = 32'b11110111011011110111111011111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011110101000000100100111101;
		b = 32'b11001111001111111010001111000111;
		correct = 32'b11001111111111111010101111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100101011110111111110011011000;
		b = 32'b10001011101010011001111111001010;
		correct = 32'b11101111111110111111111111011010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101110010100101101000101110001;
		b = 32'b00101100101001001000101111000011;
		correct = 32'b11101110111101101101101111110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100000000001100001101001110101;
		b = 32'b11011011001010011110000101101101;
		correct = 32'b11111011001011111111101101111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001011110101001010001101001000;
		b = 32'b00011011010001010001000110001001;
		correct = 32'b00011011110101011011001111001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010010111010000001001101101111;
		b = 32'b11010000001111110011000100101000;
		correct = 32'b11010010111111110011001101101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000111100101101110101111111110;
		b = 32'b10111011111111100100101010100101;
		correct = 32'b11111111111111101110101111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010000011010010001001111111100;
		b = 32'b11110111011001011100000011001011;
		correct = 32'b11110111011011011101001111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101100100011001111010110010001;
		b = 32'b00110001010010001001001110001100;
		correct = 32'b11111101110011001111011110011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00011110000011000100001001101111;
		b = 32'b01111010000100000000001100011100;
		correct = 32'b01111110000111000100001101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10000110001001111010110110110011;
		b = 32'b11001101000010001011010111000111;
		correct = 32'b11001111001011111011110111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00000010000101110100100111101011;
		b = 32'b01100101010000011010011010010010;
		correct = 32'b01100111010101111110111111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011111111111010110000101000001;
		b = 32'b00000010100101011101110010001110;
		correct = 32'b10011111111111011111110111001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111011100011010010010110010101;
		b = 32'b00011010000011101101110101101111;
		correct = 32'b10111011100011111111110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00001111100010111101101001100011;
		b = 32'b11101111010001010010111010111011;
		correct = 32'b11101111110011111111111011111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11100111000001011110111010110101;
		b = 32'b10110011100000111010111011000111;
		correct = 32'b11110111100001111110111011110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010100001101111101101100010000;
		b = 32'b10011111101110010101111101001101;
		correct = 32'b10011111101111111101111101011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011110010001001000101001110010;
		b = 32'b01011101011100001011001010101010;
		correct = 32'b11011111011101001011101011111010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101101001110100000111111010111;
		b = 32'b10001100101001010100100000100011;
		correct = 32'b11101101101111110100111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001101101000101111001000001011;
		b = 32'b10001111001111111101001110010110;
		correct = 32'b10001111101111111111001110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110101001111110000100000011110;
		b = 32'b01000111001110111001110111101001;
		correct = 32'b11110111001111111001110111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010110111010101010000110101110;
		b = 32'b11011111100010001011111001111011;
		correct = 32'b11011111111010101011111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001111110010001010011001100;
		b = 32'b11110101101111110000110101000100;
		correct = 32'b11111101111111110001110111001100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10010101010110111001000100111110;
		b = 32'b10001010000111100010111011001001;
		correct = 32'b10011111010111111011111111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001011111000111001111100011010;
		b = 32'b01001101010100100111000000100011;
		correct = 32'b01001111111100111111111100111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100110101101011011100101010;
		b = 32'b11111111000000001111001100010101;
		correct = 32'b11111111110101101111011100111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110111101101100110000010111001;
		b = 32'b00101010111010001111001001001111;
		correct = 32'b10111111111111101111001011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111101101000000100001110010101;
		b = 32'b01110100101010110111111111100110;
		correct = 32'b11111101101010110111111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010001000001011110000100101001;
		b = 32'b11000001111001001110001010100101;
		correct = 32'b11010001111001011110001110101101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11010100011110011000011010001010;
		b = 32'b01101010010000101101001011010101;
		correct = 32'b11111110011110111101011011011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101001011101010000001111101010;
		b = 32'b01010011000101010101011111010011;
		correct = 32'b11111011011101010101011111111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10011100111010111111101110010100;
		b = 32'b01010010000101100010011010011010;
		correct = 32'b11011110111111111111111110011110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101001010011010010000101000000;
		b = 32'b01110000110010101110010010101001;
		correct = 32'b01111001110011111110010111101001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000100000011011010001010000;
		b = 32'b00111010100011001101010110001111;
		correct = 32'b10111010100011011111010111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111001101100110000101101001100;
		b = 32'b00000110011101010100011101100100;
		correct = 32'b01111111111101110100111101101100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001111001111010010010001110;
		b = 32'b00011111001101100000010100001010;
		correct = 32'b00011111111101111010010110001110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000110110100001101010101100100;
		b = 32'b01010000011000001101000101000100;
		correct = 32'b11010110111100001101010101100100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011110001001100110100110001;
		b = 32'b10010011010100001001001010100011;
		correct = 32'b10111011110101001101111110110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101110010001010101000000010011;
		b = 32'b00111010000000010000010111110100;
		correct = 32'b01111110010001010101010111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01100100001010111010101011111010;
		b = 32'b01110101111111011000100111110101;
		correct = 32'b01110101111111111010101111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00101011100001000010000011000000;
		b = 32'b00010010001000111001100011000100;
		correct = 32'b00111011101001111011100011000100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011001011001010100110100110011;
		b = 32'b10001100000011100000111010011011;
		correct = 32'b11011101011011110100111110111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11101101111011100000110011011000;
		b = 32'b11110000101101000000001101000100;
		correct = 32'b11111101111111100000111111011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001111001111110001000110011101;
		b = 32'b10010111011111011000000010011010;
		correct = 32'b11011111011111111001000110011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10100000111101000111011010110001;
		b = 32'b00100111100101100011000011101110;
		correct = 32'b10100111111101100111011011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11001011000000001110100110000110;
		b = 32'b10111111101100110011010011100100;
		correct = 32'b11111111101100111111110111100110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100111001111001111110111110;
		b = 32'b10101100100111011010001110010110;
		correct = 32'b11101100111111111011111110111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10111001111101111111110110110101;
		b = 32'b10010110000111110011010110001100;
		correct = 32'b10111111111111111111110110111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010111010111111110010010100;
		b = 32'b11101110101010000111110100001100;
		correct = 32'b11101110111010111111110110011100;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100000100010010101111000001;
		b = 32'b00000100111011011000101001001001;
		correct = 32'b11011100111111011010101111001001;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111011101101111111111100111010;
		b = 32'b10000010001110101001100011101110;
		correct = 32'b11111011101111111111111111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001000010101000010000100111;
		b = 32'b01111011110110010101000111111101;
		correct = 32'b11111011110110111101010111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01011010010011011011100110000001;
		b = 32'b00000011001010100000110000001010;
		correct = 32'b01011011011011111011110110001011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101100000100111000001111101111;
		b = 32'b01010001111100001101000000011100;
		correct = 32'b11111101111100111101001111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001100101111101010011010111000;
		b = 32'b11000110001001000010010011010111;
		correct = 32'b11001110101111101010011011111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01001110011110101101001011111000;
		b = 32'b11101011011111011101000011111101;
		correct = 32'b11101111011111111101001011111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01000000001010010011111110111010;
		b = 32'b00101101110010110010000001101100;
		correct = 32'b01101101111010110011111111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111001001000000011110010011;
		b = 32'b10001001101100111001000100110010;
		correct = 32'b10101111101101111001011110110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10101111111100001101000111110110;
		b = 32'b10111101100010011001111001110001;
		correct = 32'b10111111111110011101111111110111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011111011001101011111000010000;
		b = 32'b01101000010000000101101010101000;
		correct = 32'b11111111011001101111111010111000;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010001111100000001110000001010;
		b = 32'b00011101101101010011100011001101;
		correct = 32'b00011101111101010011110011001111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11011100001001011111110111111000;
		b = 32'b10101101010011111001111001010110;
		correct = 32'b11111101011011111111111111111110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01111111111101110000100001101101;
		b = 32'b01111100110101110001011011101011;
		correct = 32'b01111111111101110001111011101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111100101010001101001110001001;
		b = 32'b11001010001101110011010111110111;
		correct = 32'b11111110101111111111011111111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01010110110010110101101100011011;
		b = 32'b11000100010100011011101101111110;
		correct = 32'b11010110110110111111101101111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000101111110110001101010111101;
		b = 32'b00101011011010001000101000111110;
		correct = 32'b11101111111110111001101010111111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11000011000101111011011010010011;
		b = 32'b11011010111111010000100101011101;
		correct = 32'b11011011111111111011111111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111010011100101001111001001000;
		b = 32'b10110110110010000111011001101111;
		correct = 32'b11111110111110101111111001101111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001010110110110011101110011101;
		b = 32'b01001100010001100110100000010000;
		correct = 32'b11001110110111110111101110011101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b01101010110101100001110101110010;
		b = 32'b11011101101111110010010101010011;
		correct = 32'b11111111111111110011110101110011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11110110101010011011011001110101;
		b = 32'b10110111110100100011001001001100;
		correct = 32'b11110111111110111011011001111101;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b11111001011101100101000010111011;
		b = 32'b00101111010100100001101001101000;
		correct = 32'b11111111011101100101101011111011;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10001000100000110101101111011101;
		b = 32'b01000101111110000001010101011010;
		correct = 32'b11001101111110110101111111011111;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b00010101101011100100110010101010;
		b = 32'b01011000001111010100001100000100;
		correct = 32'b01011101101111110100111110101110;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		a = 32'b10110000011101111010000011001010;
		b = 32'b11101011110111010110111111100000;
		correct = 32'b11111011111111111110111111101010;
			
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
		$display ("Done.");
		$finish;
	end

endmodule
